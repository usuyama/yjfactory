library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;


entity PROM is
  
  port (
    clka  : in  std_logic;
--    wea   : in  std_logic_vector(0 downto 0);
    addra : in  std_logic_vector(31 downto 0);
--    dina  : in  std_logic_vector(31 downto 0);
    douta : out std_logic_vector(31 downto 0));

end PROM;

architecture R_rom of PROM is
type rom_type is array (0 to 34) of std_logic_vector(31 downto 0);
constant rom : rom_type:=(
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00110000011000000000000000000011",--beq r0 r3 -3       9
--"10101000011000110000000000000001",--subi r3 r3 1       8
--"10000100001000100001000000000000",--add r1 r2 r2       7
--"10000100001000100000100000000000",--add r1 r2 r1       6
--"10100100000000110000000000000101",--addi r0 r3 2       5
--"10100100000000100000000000000001",--addi r0 r2 1       4
--"10100100000000010000000000000001",--addi r0 r1 1       3
--"10100100000000010000000000000001",--addi r0 r1 1       2
--"10100100000000010000000000000001"--addi r0 r1 1        1
0=>"11001011110111100000000000000011",
1=>"11001011111111110000000000000000",
2=>"11001000000111010010011100010000",
3=>"11001000000000010000000000000010",
4=>"00111111111111100000000000000000",
5=>"10100111110111100000000000000001",
6=>"01011000000000000000000000001010",
7=>"10101011110111100000000000000001",
8=>"00111011111111100000000000000000",
9=>"11000000000000000000000000000000",
10=>"11001000000000100000000000000001",
11=>"00110000001000100000000000000010",
12=>"01001111111000000000000000000000",
13=>"11001000010000000000000000000001",
14=>"10001000010000010001000000000000",
15=>"00111100001111100000000000000000",
16=>"10000100001000000001000000000000", 
17=>"00111111111111100000000000000001",
18=>"10100111110111100000000000000010",
19=>"01011000000000000000000000001010",
20=>"10101011110111100000000000000010",
21=>"00111011111111100000000000000001",
22=>"11001000000000100000000000000010",
23=>"00111000011111100000000000000000",
24=>"10001000010000110001000000000000",
25=>"00111100001111100000000000000001", 
26=>"10000100001000000001000000000000",
27=>"00111111111111100000000000000010",
28=>"10100111110111100000000000000011",
29=>"01011000000000000000000000001010",
30=>"10101011110111100000000000000011",
31=>"00111011111111100000000000000010",
32=>"00111000010111100000000000000001",
33=>"10000100001000100000100000000000",
34=>"01001111111000000000000000000000"
--"00000000000000000000000000000000",
--"10100100001000010000000000001010",
--"00111100001000010000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00111000001000100000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000"
);

signal shortened : std_logic_vector(5 downto 0):=(others=>'0');
  
begin  -- R_rom
  shortened<=addra(5 downto 0);
    douta<=rom(conv_integer(shortened));
end R_rom;
