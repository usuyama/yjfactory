library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;


entity PROM is

  port (
    clka  : in  std_logic;
--    wea   : in  std_logic_vector(0 downto 0);
    addra : in  std_logic_vector(6 downto 0);
--    dina  : in  std_logic_vector(31 downto 0);
    douta : out std_logic_vector(31 downto 0));

end PROM;

architecture R_rom of PROM is

type rom_type is array (0 to 5) of std_logic_vector(31 downto 0);
  constant rom : rom_type:=(
"11001100000111100000000000000000",
"10100100000111110000000000001111",
"11001100000111011100001101010000",
"11001100000000010000000000000100",
"11001100000000100000000000000011",
"11001100000000110000000000000010",
"11001100000001000000000000000001",
"00111111111111100000000000000000",
"10100111110111100000000000000001",
"01011000000000000000000000111001",
"10101011110111100000000000000001",
"00111011110111110000000000000000",
"11001100000000101111111000000011",
"11001000000000101111111111111111",
"01010100000000000000000000110100",
"11111100000000000000000000000000",
"11001100000000110000000000001010",
"00110000011000010000000000000110",
"11001100000000110000000000001010",
"10001000001000110000100000000000",
"11001100000000110000000000000001",
"10000100010000110001000000000000",
"01010100000000000000000000010000",
"10000100000000100000100000000000",
"01001111111000000000000000000000",
"11001100000000100000000000000000",
"01010100000000000000000000010000",
"11001100000000100000000000001010",
"00110000010000010000000000010101",
"00111100001111100000000000000000",
"00111111111111100000000000000001",
"10100111110111100000000000000010",
"01011000000000000000000000011001",
"10101011110111100000000000000010",
"00111011110111110000000000000001",
"00111100001111100000000000000001",
"00111111111111100000000000000010",
"10100111110111100000000000000011",
"01011000000000000000000000011011",
"10101011110111100000000000000011",
"00111011110111110000000000000010",
"11001100000000010000000000001010",
"00111011110000100000000000000001",
"10001100010000010000100000000000",
"00111011110000100000000000000000",
"10001000010000010000100000000000",
"11001100000000100000000000110000",
"10000100001000100000100000000000",
"01010100000000000000000010011100",
"11001100000000100000000000110000",
"10000100001000100000100000000000",
"01010100000000000000000010011100",
"00101000001000100000000000000011",
"11001100000000010000000000000001",
"01010100000000000000000000011011",
"11001100000000010000000000000000",
"01010100000000000000000000011011",
"10000100001000100010100000000000",
"10000100001000110011000000000000",
"10000100001001000011100000000000",
"10000100010000110100000000000000",
"10000100010001000100100000000000",
"10000100011001000101000000000000",
"10000100101001100101100000000000",
"10000100101001110110000000000000",
"10000100101010000110100000000000",
"10000100101010010111000000000000",
"10000100101010100111100000000000",
"10000100110001111000000000000000",
"10000100110010001000100000000000",
"10000100110010011001000000000000",
"10000100110010101001100000000000",
"10000100111010001010000000000000",
"10000100111010011010100000000000",
"10000100111010101011000000000000",
"10000101000010011011100000000000",
"10000101000010101100000000000000",
"10000101001010101100100000000000",
"10000101011011001101000000000000",
"10000101011011011101100000000000",
"00111111011111100000000000000000",
"10000101011011101101100000000000",
"00111111011111100000000000000001",
"10000101011011111101100000000000",
"00111111011111100000000000000010",
"10000101011100001101100000000000",
"00111111011111100000000000000011",
"10000101011100011101100000000000",
"00111111011111100000000000000100",
"10000101011100101101100000000000",
"00111111011111100000000000000101",
"10000101011100111101100000000000",
"00111111011111100000000000000110",
"10000101011101001101100000000000",
"00111111011111100000000000000111",
"10000101011101011101100000000000",
"00111111011111100000000000001000",
"10000101011101101101100000000000",
"00111111011111100000000000001001",
"10000101011101111101100000000000",
"00111111011111100000000000001010",
"10000101011110001101100000000000",
"00111111011111100000000000001011",
"10000101011110011101100000000000",
"10000100001000100000100000000000",
"10000100001000110000100000000000",
"10000100001001000000100000000000",
"10000100001001010000100000000000",
"10000100001001100000100000000000",
"10000100001001110000100000000000",
"10000100001010000000100000000000",
"10000100001010010000100000000000",
"10000100001010100000100000000000",
"10000100001010110000100000000000",
"10000100001011000000100000000000",
"10000100001011010000100000000000",
"10000100001011100000100000000000",
"10000100001011110000100000000000",
"10000100001100000000100000000000",
"10000100001100010000100000000000",
"10000100001100100000100000000000",
"10000100001100110000100000000000",
"10000100001101000000100000000000",
"10000100001101010000100000000000",
"10000100001101100000100000000000",
"10000100001101110000100000000000",
"10000100001110000000100000000000",
"10000100001110010000100000000000",
"10000100001110100000100000000000",
"00111011110000100000000000000000",
"10000100001000100000100000000000",
"00111011110000100000000000000001",
"10000100001000100000100000000000",
"00111011110000100000000000000010",
"10000100001000100000100000000000",
"00111011110000100000000000000011",
"10000100001000100000100000000000",
"00111011110000100000000000000100",
"10000100001000100000100000000000",
"00111011110000100000000000000101",
"10000100001000100000100000000000",
"00111011110000100000000000000110",
"10000100001000100000100000000000",
"00111011110000100000000000000111",
"10000100001000100000100000000000",
"00111011110000100000000000001000",
"10000100001000100000100000000000",
"00111011110000100000000000001001",
"10000100001000100000100000000000",
"00111011110000100000000000001010",
"10000100001000100000100000000000",
"00111011110000100000000000001011",
"10000100001000100000100000000000",
"10000100001110110000100000000000",
"10001000000000010000100000000000",
"01001111111000000000000000000000",
"11010000001000000000000000000000",
"01001111111000000000000000000000",
"11001100000000110000000000000000",
"10000111101000110010000000000000",
"00111100010001000000000000000000",
"10100100011000110000000000000001",
"00110000001000111111111111111101",
"10000100000111010000100000000000",
"10000111101000111110100000000000",
"01001111111000000000000000000000",
"11001100000000110000000000000000",
"10000111101000110010000000000000",
"10110000000001000000000000000000",
"10100100011000110000000000000001",
"00110000001000111111111111111101",
"10000100000111010000100000000000",
"10000111101000111110100000000000",
"01001111111000000000000000000000",
"01100000001000000000000000000000",
"01001111111000000000000000000000",
"01100100000000010000000000000000",
"01001111111000000000000000000000",
"11110000000000000000000000000000",
"01001111111000000000000000000000",
"11110100000000000000000000000000",
"01001111111000000000000000000000",
"11001100000000010000000000000000",
"11001100000000100000000000000000",
"11000100000000010000000000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001111111000000000000000000000",
"11001100000000010000000000000000",
"11001100000000100000000000000000",
"11000100000000010000000000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01111100001000000000000000000000",
"01001111111000000000000000000000",
"11111000000000000000000000000000",
"01001111111000000000000000000000",
"00011000000000000000000000000000",
"01001111111000000000000000000000"
	-- entry:                
);                               
signal read_a : std_logic_vector(6 downto 0);
signal shortened : std_logic_vector(6 downto 0):=(others=>'0');
begin  -- R_rom
  process(clk)
    if (clk'event and clk='1')then
      read_a<=addra;
    end if;
  end process;
  shortened<=read_a(6 downto 0);
    douta<=rom(conv_integer(shortened));
end R_rom;






