library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;


entity PROM is

  port (
    clka  : in  std_logic;
--    wea   : in  std_logic_vector(0 downto 0);
    addra : in  std_logic_vector(6 downto 0);
--    dina  : in  std_logic_vector(31 downto 0);
    douta : out std_logic_vector(31 downto 0));

end PROM;

architecture R_rom of PROM is

type rom_type is array (0 to 10832) of std_logic_vector(31 downto 0);
  constant rom : rom_type:=(
	-- entry:
"00000000000000000000000000000000",	-- 0: 	nop
"11001100000111100000000000000000",	-- 1: 	lli	%sp, 0
"10100100000111110000001111110100",	-- 2: 	addi	%ra, %r0, halt
"11001100000111011100001101010000",	-- 3: 	lli	%hp, 50000
"11001100000000010000000000000001",	-- 4: 	lli	%r1, 1
"11001100000000100000000000000000",	-- 5: 	lli	%r2, 0
"00111111111111100000000000000000",	-- 6: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 7: 	addi	%sp, %sp, 1
"01011000000000000010101000011010",	-- 8: 	jal	yj_create_array
"10101011110111100000000000000001",	-- 9: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 10: 	lw	%ra, [%sp + 0]
"11001100000000100000000000000000",	-- 11: 	lli	%r2, 0
"00010100000000000000000000000000",	-- 12: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 13: 	lhif	%f0, 0.000000
"00111100001111100000000000000000",	-- 14: 	sw	%r1, [%sp + 0]
"10000100000000100000100000000000",	-- 15: 	add	%r1, %r0, %r2
"00111111111111100000000000000001",	-- 16: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 17: 	addi	%sp, %sp, 2
"01011000000000000010101000100010",	-- 18: 	jal	yj_create_float_array
"10101011110111100000000000000010",	-- 19: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 20: 	lw	%ra, [%sp + 1]
"11001100000000100000000000111100",	-- 21: 	lli	%r2, 60
"11001100000000110000000000000000",	-- 22: 	lli	%r3, 0
"11001100000001000000000000000000",	-- 23: 	lli	%r4, 0
"11001100000001010000000000000000",	-- 24: 	lli	%r5, 0
"11001100000001100000000000000000",	-- 25: 	lli	%r6, 0
"11001100000001110000000000000000",	-- 26: 	lli	%r7, 0
"10000100000111010100000000000000",	-- 27: 	add	%r8, %r0, %hp
"10100111101111010000000000001011",	-- 28: 	addi	%hp, %hp, 11
"00111100001010000000000000001010",	-- 29: 	sw	%r1, [%r8 + 10]
"00111100001010000000000000001001",	-- 30: 	sw	%r1, [%r8 + 9]
"00111100001010000000000000001000",	-- 31: 	sw	%r1, [%r8 + 8]
"00111100001010000000000000000111",	-- 32: 	sw	%r1, [%r8 + 7]
"00111100111010000000000000000110",	-- 33: 	sw	%r7, [%r8 + 6]
"00111100001010000000000000000101",	-- 34: 	sw	%r1, [%r8 + 5]
"00111100001010000000000000000100",	-- 35: 	sw	%r1, [%r8 + 4]
"00111100110010000000000000000011",	-- 36: 	sw	%r6, [%r8 + 3]
"00111100101010000000000000000010",	-- 37: 	sw	%r5, [%r8 + 2]
"00111100100010000000000000000001",	-- 38: 	sw	%r4, [%r8 + 1]
"00111100011010000000000000000000",	-- 39: 	sw	%r3, [%r8 + 0]
"10000100000010000000100000000000",	-- 40: 	add	%r1, %r0, %r8
"10000100000000101101000000000000",	-- 41: 	add	%r26, %r0, %r2
"10000100000000010001000000000000",	-- 42: 	add	%r2, %r0, %r1
"10000100000110100000100000000000",	-- 43: 	add	%r1, %r0, %r26
"00111111111111100000000000000001",	-- 44: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 45: 	addi	%sp, %sp, 2
"01011000000000000010101000011010",	-- 46: 	jal	yj_create_array
"10101011110111100000000000000010",	-- 47: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 48: 	lw	%ra, [%sp + 1]
"11001100000000100000000000000011",	-- 49: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 50: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 51: 	lhif	%f0, 0.000000
"00111100001111100000000000000001",	-- 52: 	sw	%r1, [%sp + 1]
"10000100000000100000100000000000",	-- 53: 	add	%r1, %r0, %r2
"00111111111111100000000000000010",	-- 54: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 55: 	addi	%sp, %sp, 3
"01011000000000000010101000100010",	-- 56: 	jal	yj_create_float_array
"10101011110111100000000000000011",	-- 57: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 58: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000011",	-- 59: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 60: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 61: 	lhif	%f0, 0.000000
"00111100001111100000000000000010",	-- 62: 	sw	%r1, [%sp + 2]
"10000100000000100000100000000000",	-- 63: 	add	%r1, %r0, %r2
"00111111111111100000000000000011",	-- 64: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 65: 	addi	%sp, %sp, 4
"01011000000000000010101000100010",	-- 66: 	jal	yj_create_float_array
"10101011110111100000000000000100",	-- 67: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 68: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000011",	-- 69: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 70: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 71: 	lhif	%f0, 0.000000
"00111100001111100000000000000011",	-- 72: 	sw	%r1, [%sp + 3]
"10000100000000100000100000000000",	-- 73: 	add	%r1, %r0, %r2
"00111111111111100000000000000100",	-- 74: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 75: 	addi	%sp, %sp, 5
"01011000000000000010101000100010",	-- 76: 	jal	yj_create_float_array
"10101011110111100000000000000101",	-- 77: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 78: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000001",	-- 79: 	lli	%r2, 1
"00010100000000000000000000000000",	-- 80: 	llif	%f0, 255.000000
"00010000000000000100001101111111",	-- 81: 	lhif	%f0, 255.000000
"00111100001111100000000000000100",	-- 82: 	sw	%r1, [%sp + 4]
"10000100000000100000100000000000",	-- 83: 	add	%r1, %r0, %r2
"00111111111111100000000000000101",	-- 84: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 85: 	addi	%sp, %sp, 6
"01011000000000000010101000100010",	-- 86: 	jal	yj_create_float_array
"10101011110111100000000000000110",	-- 87: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 88: 	lw	%ra, [%sp + 5]
"11001100000000100000000000110010",	-- 89: 	lli	%r2, 50
"11001100000000110000000000000001",	-- 90: 	lli	%r3, 1
"11001100000001001111111111111111",	-- 91: 	lli	%r4, -1
"11001000000001001111111111111111",	-- 92: 	lhi	%r4, -1
"00111100001111100000000000000101",	-- 93: 	sw	%r1, [%sp + 5]
"00111100010111100000000000000110",	-- 94: 	sw	%r2, [%sp + 6]
"10000100000001000001000000000000",	-- 95: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 96: 	add	%r1, %r0, %r3
"00111111111111100000000000000111",	-- 97: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 98: 	addi	%sp, %sp, 8
"01011000000000000010101000011010",	-- 99: 	jal	yj_create_array
"10101011110111100000000000001000",	-- 100: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 101: 	lw	%ra, [%sp + 7]
"10000100000000010001000000000000",	-- 102: 	add	%r2, %r0, %r1
"00111011110000010000000000000110",	-- 103: 	lw	%r1, [%sp + 6]
"00111111111111100000000000000111",	-- 104: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 105: 	addi	%sp, %sp, 8
"01011000000000000010101000011010",	-- 106: 	jal	yj_create_array
"10101011110111100000000000001000",	-- 107: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 108: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000001",	-- 109: 	lli	%r2, 1
"11001100000000110000000000000001",	-- 110: 	lli	%r3, 1
"11001100000001000000000000000000",	-- 111: 	lli	%r4, 0
"10000100001001000010000000000000",	-- 112: 	add	%r4, %r1, %r4
"00111000100001000000000000000000",	-- 113: 	lw	%r4, [%r4 + 0]
"00111100001111100000000000000111",	-- 114: 	sw	%r1, [%sp + 7]
"00111100010111100000000000001000",	-- 115: 	sw	%r2, [%sp + 8]
"10000100000001000001000000000000",	-- 116: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 117: 	add	%r1, %r0, %r3
"00111111111111100000000000001001",	-- 118: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 119: 	addi	%sp, %sp, 10
"01011000000000000010101000011010",	-- 120: 	jal	yj_create_array
"10101011110111100000000000001010",	-- 121: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 122: 	lw	%ra, [%sp + 9]
"10000100000000010001000000000000",	-- 123: 	add	%r2, %r0, %r1
"00111011110000010000000000001000",	-- 124: 	lw	%r1, [%sp + 8]
"00111111111111100000000000001001",	-- 125: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 126: 	addi	%sp, %sp, 10
"01011000000000000010101000011010",	-- 127: 	jal	yj_create_array
"10101011110111100000000000001010",	-- 128: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 129: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000001",	-- 130: 	lli	%r2, 1
"00010100000000000000000000000000",	-- 131: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 132: 	lhif	%f0, 0.000000
"00111100001111100000000000001001",	-- 133: 	sw	%r1, [%sp + 9]
"10000100000000100000100000000000",	-- 134: 	add	%r1, %r0, %r2
"00111111111111100000000000001010",	-- 135: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 136: 	addi	%sp, %sp, 11
"01011000000000000010101000100010",	-- 137: 	jal	yj_create_float_array
"10101011110111100000000000001011",	-- 138: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 139: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000001",	-- 140: 	lli	%r2, 1
"11001100000000110000000000000000",	-- 141: 	lli	%r3, 0
"00111100001111100000000000001010",	-- 142: 	sw	%r1, [%sp + 10]
"10000100000000100000100000000000",	-- 143: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 144: 	add	%r2, %r0, %r3
"00111111111111100000000000001011",	-- 145: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 146: 	addi	%sp, %sp, 12
"01011000000000000010101000011010",	-- 147: 	jal	yj_create_array
"10101011110111100000000000001100",	-- 148: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 149: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000001",	-- 150: 	lli	%r2, 1
"00010100000000000110101100101000",	-- 151: 	llif	%f0, 1000000000.000000
"00010000000000000100111001101110",	-- 152: 	lhif	%f0, 1000000000.000000
"00111100001111100000000000001011",	-- 153: 	sw	%r1, [%sp + 11]
"10000100000000100000100000000000",	-- 154: 	add	%r1, %r0, %r2
"00111111111111100000000000001100",	-- 155: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 156: 	addi	%sp, %sp, 13
"01011000000000000010101000100010",	-- 157: 	jal	yj_create_float_array
"10101011110111100000000000001101",	-- 158: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 159: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000011",	-- 160: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 161: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 162: 	lhif	%f0, 0.000000
"00111100001111100000000000001100",	-- 163: 	sw	%r1, [%sp + 12]
"10000100000000100000100000000000",	-- 164: 	add	%r1, %r0, %r2
"00111111111111100000000000001101",	-- 165: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 166: 	addi	%sp, %sp, 14
"01011000000000000010101000100010",	-- 167: 	jal	yj_create_float_array
"10101011110111100000000000001110",	-- 168: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 169: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000001",	-- 170: 	lli	%r2, 1
"11001100000000110000000000000000",	-- 171: 	lli	%r3, 0
"00111100001111100000000000001101",	-- 172: 	sw	%r1, [%sp + 13]
"10000100000000100000100000000000",	-- 173: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 174: 	add	%r2, %r0, %r3
"00111111111111100000000000001110",	-- 175: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 176: 	addi	%sp, %sp, 15
"01011000000000000010101000011010",	-- 177: 	jal	yj_create_array
"10101011110111100000000000001111",	-- 178: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 179: 	lw	%ra, [%sp + 14]
"11001100000000100000000000000011",	-- 180: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 181: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 182: 	lhif	%f0, 0.000000
"00111100001111100000000000001110",	-- 183: 	sw	%r1, [%sp + 14]
"10000100000000100000100000000000",	-- 184: 	add	%r1, %r0, %r2
"00111111111111100000000000001111",	-- 185: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 186: 	addi	%sp, %sp, 16
"01011000000000000010101000100010",	-- 187: 	jal	yj_create_float_array
"10101011110111100000000000010000",	-- 188: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 189: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000011",	-- 190: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 191: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 192: 	lhif	%f0, 0.000000
"00111100001111100000000000001111",	-- 193: 	sw	%r1, [%sp + 15]
"10000100000000100000100000000000",	-- 194: 	add	%r1, %r0, %r2
"00111111111111100000000000010000",	-- 195: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 196: 	addi	%sp, %sp, 17
"01011000000000000010101000100010",	-- 197: 	jal	yj_create_float_array
"10101011110111100000000000010001",	-- 198: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 199: 	lw	%ra, [%sp + 16]
"11001100000000100000000000000011",	-- 200: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 201: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 202: 	lhif	%f0, 0.000000
"00111100001111100000000000010000",	-- 203: 	sw	%r1, [%sp + 16]
"10000100000000100000100000000000",	-- 204: 	add	%r1, %r0, %r2
"00111111111111100000000000010001",	-- 205: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 206: 	addi	%sp, %sp, 18
"01011000000000000010101000100010",	-- 207: 	jal	yj_create_float_array
"10101011110111100000000000010010",	-- 208: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 209: 	lw	%ra, [%sp + 17]
"11001100000000100000000000000011",	-- 210: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 211: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 212: 	lhif	%f0, 0.000000
"00111100001111100000000000010001",	-- 213: 	sw	%r1, [%sp + 17]
"10000100000000100000100000000000",	-- 214: 	add	%r1, %r0, %r2
"00111111111111100000000000010010",	-- 215: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 216: 	addi	%sp, %sp, 19
"01011000000000000010101000100010",	-- 217: 	jal	yj_create_float_array
"10101011110111100000000000010011",	-- 218: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 219: 	lw	%ra, [%sp + 18]
"11001100000000100000000000000010",	-- 220: 	lli	%r2, 2
"11001100000000110000000000000000",	-- 221: 	lli	%r3, 0
"00111100001111100000000000010010",	-- 222: 	sw	%r1, [%sp + 18]
"10000100000000100000100000000000",	-- 223: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 224: 	add	%r2, %r0, %r3
"00111111111111100000000000010011",	-- 225: 	sw	%ra, [%sp + 19]
"10100111110111100000000000010100",	-- 226: 	addi	%sp, %sp, 20
"01011000000000000010101000011010",	-- 227: 	jal	yj_create_array
"10101011110111100000000000010100",	-- 228: 	subi	%sp, %sp, 20
"00111011110111110000000000010011",	-- 229: 	lw	%ra, [%sp + 19]
"11001100000000100000000000000010",	-- 230: 	lli	%r2, 2
"11001100000000110000000000000000",	-- 231: 	lli	%r3, 0
"00111100001111100000000000010011",	-- 232: 	sw	%r1, [%sp + 19]
"10000100000000100000100000000000",	-- 233: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 234: 	add	%r2, %r0, %r3
"00111111111111100000000000010100",	-- 235: 	sw	%ra, [%sp + 20]
"10100111110111100000000000010101",	-- 236: 	addi	%sp, %sp, 21
"01011000000000000010101000011010",	-- 237: 	jal	yj_create_array
"10101011110111100000000000010101",	-- 238: 	subi	%sp, %sp, 21
"00111011110111110000000000010100",	-- 239: 	lw	%ra, [%sp + 20]
"11001100000000100000000000000001",	-- 240: 	lli	%r2, 1
"00010100000000000000000000000000",	-- 241: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 242: 	lhif	%f0, 0.000000
"00111100001111100000000000010100",	-- 243: 	sw	%r1, [%sp + 20]
"10000100000000100000100000000000",	-- 244: 	add	%r1, %r0, %r2
"00111111111111100000000000010101",	-- 245: 	sw	%ra, [%sp + 21]
"10100111110111100000000000010110",	-- 246: 	addi	%sp, %sp, 22
"01011000000000000010101000100010",	-- 247: 	jal	yj_create_float_array
"10101011110111100000000000010110",	-- 248: 	subi	%sp, %sp, 22
"00111011110111110000000000010101",	-- 249: 	lw	%ra, [%sp + 21]
"11001100000000100000000000000011",	-- 250: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 251: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 252: 	lhif	%f0, 0.000000
"00111100001111100000000000010101",	-- 253: 	sw	%r1, [%sp + 21]
"10000100000000100000100000000000",	-- 254: 	add	%r1, %r0, %r2
"00111111111111100000000000010110",	-- 255: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 256: 	addi	%sp, %sp, 23
"01011000000000000010101000100010",	-- 257: 	jal	yj_create_float_array
"10101011110111100000000000010111",	-- 258: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 259: 	lw	%ra, [%sp + 22]
"11001100000000100000000000000011",	-- 260: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 261: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 262: 	lhif	%f0, 0.000000
"00111100001111100000000000010110",	-- 263: 	sw	%r1, [%sp + 22]
"10000100000000100000100000000000",	-- 264: 	add	%r1, %r0, %r2
"00111111111111100000000000010111",	-- 265: 	sw	%ra, [%sp + 23]
"10100111110111100000000000011000",	-- 266: 	addi	%sp, %sp, 24
"01011000000000000010101000100010",	-- 267: 	jal	yj_create_float_array
"10101011110111100000000000011000",	-- 268: 	subi	%sp, %sp, 24
"00111011110111110000000000010111",	-- 269: 	lw	%ra, [%sp + 23]
"11001100000000100000000000000011",	-- 270: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 271: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 272: 	lhif	%f0, 0.000000
"00111100001111100000000000010111",	-- 273: 	sw	%r1, [%sp + 23]
"10000100000000100000100000000000",	-- 274: 	add	%r1, %r0, %r2
"00111111111111100000000000011000",	-- 275: 	sw	%ra, [%sp + 24]
"10100111110111100000000000011001",	-- 276: 	addi	%sp, %sp, 25
"01011000000000000010101000100010",	-- 277: 	jal	yj_create_float_array
"10101011110111100000000000011001",	-- 278: 	subi	%sp, %sp, 25
"00111011110111110000000000011000",	-- 279: 	lw	%ra, [%sp + 24]
"11001100000000100000000000000011",	-- 280: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 281: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 282: 	lhif	%f0, 0.000000
"00111100001111100000000000011000",	-- 283: 	sw	%r1, [%sp + 24]
"10000100000000100000100000000000",	-- 284: 	add	%r1, %r0, %r2
"00111111111111100000000000011001",	-- 285: 	sw	%ra, [%sp + 25]
"10100111110111100000000000011010",	-- 286: 	addi	%sp, %sp, 26
"01011000000000000010101000100010",	-- 287: 	jal	yj_create_float_array
"10101011110111100000000000011010",	-- 288: 	subi	%sp, %sp, 26
"00111011110111110000000000011001",	-- 289: 	lw	%ra, [%sp + 25]
"11001100000000100000000000000011",	-- 290: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 291: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 292: 	lhif	%f0, 0.000000
"00111100001111100000000000011001",	-- 293: 	sw	%r1, [%sp + 25]
"10000100000000100000100000000000",	-- 294: 	add	%r1, %r0, %r2
"00111111111111100000000000011010",	-- 295: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 296: 	addi	%sp, %sp, 27
"01011000000000000010101000100010",	-- 297: 	jal	yj_create_float_array
"10101011110111100000000000011011",	-- 298: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 299: 	lw	%ra, [%sp + 26]
"11001100000000100000000000000011",	-- 300: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 301: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 302: 	lhif	%f0, 0.000000
"00111100001111100000000000011010",	-- 303: 	sw	%r1, [%sp + 26]
"10000100000000100000100000000000",	-- 304: 	add	%r1, %r0, %r2
"00111111111111100000000000011011",	-- 305: 	sw	%ra, [%sp + 27]
"10100111110111100000000000011100",	-- 306: 	addi	%sp, %sp, 28
"01011000000000000010101000100010",	-- 307: 	jal	yj_create_float_array
"10101011110111100000000000011100",	-- 308: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 309: 	lw	%ra, [%sp + 27]
"11001100000000100000000000000000",	-- 310: 	lli	%r2, 0
"00010100000000000000000000000000",	-- 311: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 312: 	lhif	%f0, 0.000000
"00111100001111100000000000011011",	-- 313: 	sw	%r1, [%sp + 27]
"10000100000000100000100000000000",	-- 314: 	add	%r1, %r0, %r2
"00111111111111100000000000011100",	-- 315: 	sw	%ra, [%sp + 28]
"10100111110111100000000000011101",	-- 316: 	addi	%sp, %sp, 29
"01011000000000000010101000100010",	-- 317: 	jal	yj_create_float_array
"10101011110111100000000000011101",	-- 318: 	subi	%sp, %sp, 29
"00111011110111110000000000011100",	-- 319: 	lw	%ra, [%sp + 28]
"10000100000000010001000000000000",	-- 320: 	add	%r2, %r0, %r1
"11001100000000010000000000000000",	-- 321: 	lli	%r1, 0
"00111100010111100000000000011100",	-- 322: 	sw	%r2, [%sp + 28]
"00111111111111100000000000011101",	-- 323: 	sw	%ra, [%sp + 29]
"10100111110111100000000000011110",	-- 324: 	addi	%sp, %sp, 30
"01011000000000000010101000011010",	-- 325: 	jal	yj_create_array
"10101011110111100000000000011110",	-- 326: 	subi	%sp, %sp, 30
"00111011110111110000000000011101",	-- 327: 	lw	%ra, [%sp + 29]
"11001100000000100000000000000000",	-- 328: 	lli	%r2, 0
"10000100000111010001100000000000",	-- 329: 	add	%r3, %r0, %hp
"10100111101111010000000000000010",	-- 330: 	addi	%hp, %hp, 2
"00111100001000110000000000000001",	-- 331: 	sw	%r1, [%r3 + 1]
"00111011110000010000000000011100",	-- 332: 	lw	%r1, [%sp + 28]
"00111100001000110000000000000000",	-- 333: 	sw	%r1, [%r3 + 0]
"10000100000000110000100000000000",	-- 334: 	add	%r1, %r0, %r3
"10000100000000101101000000000000",	-- 335: 	add	%r26, %r0, %r2
"10000100000000010001000000000000",	-- 336: 	add	%r2, %r0, %r1
"10000100000110100000100000000000",	-- 337: 	add	%r1, %r0, %r26
"00111111111111100000000000011101",	-- 338: 	sw	%ra, [%sp + 29]
"10100111110111100000000000011110",	-- 339: 	addi	%sp, %sp, 30
"01011000000000000010101000011010",	-- 340: 	jal	yj_create_array
"10101011110111100000000000011110",	-- 341: 	subi	%sp, %sp, 30
"00111011110111110000000000011101",	-- 342: 	lw	%ra, [%sp + 29]
"10000100000000010001000000000000",	-- 343: 	add	%r2, %r0, %r1
"11001100000000010000000000000101",	-- 344: 	lli	%r1, 5
"00111111111111100000000000011101",	-- 345: 	sw	%ra, [%sp + 29]
"10100111110111100000000000011110",	-- 346: 	addi	%sp, %sp, 30
"01011000000000000010101000011010",	-- 347: 	jal	yj_create_array
"10101011110111100000000000011110",	-- 348: 	subi	%sp, %sp, 30
"00111011110111110000000000011101",	-- 349: 	lw	%ra, [%sp + 29]
"11001100000000100000000000000000",	-- 350: 	lli	%r2, 0
"00010100000000000000000000000000",	-- 351: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 352: 	lhif	%f0, 0.000000
"00111100001111100000000000011101",	-- 353: 	sw	%r1, [%sp + 29]
"10000100000000100000100000000000",	-- 354: 	add	%r1, %r0, %r2
"00111111111111100000000000011110",	-- 355: 	sw	%ra, [%sp + 30]
"10100111110111100000000000011111",	-- 356: 	addi	%sp, %sp, 31
"01011000000000000010101000100010",	-- 357: 	jal	yj_create_float_array
"10101011110111100000000000011111",	-- 358: 	subi	%sp, %sp, 31
"00111011110111110000000000011110",	-- 359: 	lw	%ra, [%sp + 30]
"11001100000000100000000000000011",	-- 360: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 361: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 362: 	lhif	%f0, 0.000000
"00111100001111100000000000011110",	-- 363: 	sw	%r1, [%sp + 30]
"10000100000000100000100000000000",	-- 364: 	add	%r1, %r0, %r2
"00111111111111100000000000011111",	-- 365: 	sw	%ra, [%sp + 31]
"10100111110111100000000000100000",	-- 366: 	addi	%sp, %sp, 32
"01011000000000000010101000100010",	-- 367: 	jal	yj_create_float_array
"10101011110111100000000000100000",	-- 368: 	subi	%sp, %sp, 32
"00111011110111110000000000011111",	-- 369: 	lw	%ra, [%sp + 31]
"11001100000000100000000000111100",	-- 370: 	lli	%r2, 60
"00111011110000110000000000011110",	-- 371: 	lw	%r3, [%sp + 30]
"00111100001111100000000000011111",	-- 372: 	sw	%r1, [%sp + 31]
"10000100000000100000100000000000",	-- 373: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 374: 	add	%r2, %r0, %r3
"00111111111111100000000000100000",	-- 375: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 376: 	addi	%sp, %sp, 33
"01011000000000000010101000011010",	-- 377: 	jal	yj_create_array
"10101011110111100000000000100001",	-- 378: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 379: 	lw	%ra, [%sp + 32]
"10000100000111010001000000000000",	-- 380: 	add	%r2, %r0, %hp
"10100111101111010000000000000010",	-- 381: 	addi	%hp, %hp, 2
"00111100001000100000000000000001",	-- 382: 	sw	%r1, [%r2 + 1]
"00111011110000010000000000011111",	-- 383: 	lw	%r1, [%sp + 31]
"00111100001000100000000000000000",	-- 384: 	sw	%r1, [%r2 + 0]
"10000100000000100000100000000000",	-- 385: 	add	%r1, %r0, %r2
"11001100000000100000000000000000",	-- 386: 	lli	%r2, 0
"00010100000000000000000000000000",	-- 387: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 388: 	lhif	%f0, 0.000000
"00111100001111100000000000100000",	-- 389: 	sw	%r1, [%sp + 32]
"10000100000000100000100000000000",	-- 390: 	add	%r1, %r0, %r2
"00111111111111100000000000100001",	-- 391: 	sw	%ra, [%sp + 33]
"10100111110111100000000000100010",	-- 392: 	addi	%sp, %sp, 34
"01011000000000000010101000100010",	-- 393: 	jal	yj_create_float_array
"10101011110111100000000000100010",	-- 394: 	subi	%sp, %sp, 34
"00111011110111110000000000100001",	-- 395: 	lw	%ra, [%sp + 33]
"10000100000000010001000000000000",	-- 396: 	add	%r2, %r0, %r1
"11001100000000010000000000000000",	-- 397: 	lli	%r1, 0
"00111100010111100000000000100001",	-- 398: 	sw	%r2, [%sp + 33]
"00111111111111100000000000100010",	-- 399: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 400: 	addi	%sp, %sp, 35
"01011000000000000010101000011010",	-- 401: 	jal	yj_create_array
"10101011110111100000000000100011",	-- 402: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 403: 	lw	%ra, [%sp + 34]
"10000100000111010001000000000000",	-- 404: 	add	%r2, %r0, %hp
"10100111101111010000000000000010",	-- 405: 	addi	%hp, %hp, 2
"00111100001000100000000000000001",	-- 406: 	sw	%r1, [%r2 + 1]
"00111011110000010000000000100001",	-- 407: 	lw	%r1, [%sp + 33]
"00111100001000100000000000000000",	-- 408: 	sw	%r1, [%r2 + 0]
"10000100000000100000100000000000",	-- 409: 	add	%r1, %r0, %r2
"11001100000000100000000010110100",	-- 410: 	lli	%r2, 180
"11001100000000110000000000000000",	-- 411: 	lli	%r3, 0
"00010100000000000000000000000000",	-- 412: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 413: 	lhif	%f0, 0.000000
"10000100000111010010000000000000",	-- 414: 	add	%r4, %r0, %hp
"10100111101111010000000000000011",	-- 415: 	addi	%hp, %hp, 3
"10110000000001000000000000000010",	-- 416: 	sf	%f0, [%r4 + 2]
"00111100001001000000000000000001",	-- 417: 	sw	%r1, [%r4 + 1]
"00111100011001000000000000000000",	-- 418: 	sw	%r3, [%r4 + 0]
"10000100000001000000100000000000",	-- 419: 	add	%r1, %r0, %r4
"10000100000000101101000000000000",	-- 420: 	add	%r26, %r0, %r2
"10000100000000010001000000000000",	-- 421: 	add	%r2, %r0, %r1
"10000100000110100000100000000000",	-- 422: 	add	%r1, %r0, %r26
"00111111111111100000000000100010",	-- 423: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 424: 	addi	%sp, %sp, 35
"01011000000000000010101000011010",	-- 425: 	jal	yj_create_array
"10101011110111100000000000100011",	-- 426: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 427: 	lw	%ra, [%sp + 34]
"11001100000000100000000000000001",	-- 428: 	lli	%r2, 1
"11001100000000110000000000000000",	-- 429: 	lli	%r3, 0
"00111100001111100000000000100010",	-- 430: 	sw	%r1, [%sp + 34]
"10000100000000100000100000000000",	-- 431: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 432: 	add	%r2, %r0, %r3
"00111111111111100000000000100011",	-- 433: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 434: 	addi	%sp, %sp, 36
"01011000000000000010101000011010",	-- 435: 	jal	yj_create_array
"10101011110111100000000000100100",	-- 436: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 437: 	lw	%ra, [%sp + 35]
"10000100000111010001000000000000",	-- 438: 	add	%r2, %r0, %hp
"10100111101111010000000000000110",	-- 439: 	addi	%hp, %hp, 6
"10100100000000110000011011001000",	-- 440: 	addi	%r3, %r0, read_screen_settings.2695
"00111100011000100000000000000000",	-- 441: 	sw	%r3, [%r2 + 0]
"00111011110000110000000000000011",	-- 442: 	lw	%r3, [%sp + 3]
"00111100011000100000000000000101",	-- 443: 	sw	%r3, [%r2 + 5]
"00111011110001000000000000011010",	-- 444: 	lw	%r4, [%sp + 26]
"00111100100000100000000000000100",	-- 445: 	sw	%r4, [%r2 + 4]
"00111011110001010000000000011001",	-- 446: 	lw	%r5, [%sp + 25]
"00111100101000100000000000000011",	-- 447: 	sw	%r5, [%r2 + 3]
"00111011110001100000000000011000",	-- 448: 	lw	%r6, [%sp + 24]
"00111100110000100000000000000010",	-- 449: 	sw	%r6, [%r2 + 2]
"00111011110001110000000000000010",	-- 450: 	lw	%r7, [%sp + 2]
"00111100111000100000000000000001",	-- 451: 	sw	%r7, [%r2 + 1]
"10000100000111010011100000000000",	-- 452: 	add	%r7, %r0, %hp
"10100111101111010000000000000011",	-- 453: 	addi	%hp, %hp, 3
"10100100000010000000011110011011",	-- 454: 	addi	%r8, %r0, read_light.2697
"00111101000001110000000000000000",	-- 455: 	sw	%r8, [%r7 + 0]
"00111011110010000000000000000100",	-- 456: 	lw	%r8, [%sp + 4]
"00111101000001110000000000000010",	-- 457: 	sw	%r8, [%r7 + 2]
"00111011110010010000000000000101",	-- 458: 	lw	%r9, [%sp + 5]
"00111101001001110000000000000001",	-- 459: 	sw	%r9, [%r7 + 1]
"10000100000111010101000000000000",	-- 460: 	add	%r10, %r0, %hp
"10100111101111010000000000000010",	-- 461: 	addi	%hp, %hp, 2
"10100100000010110000100100011010",	-- 462: 	addi	%r11, %r0, read_nth_object.2702
"00111101011010100000000000000000",	-- 463: 	sw	%r11, [%r10 + 0]
"00111011110010110000000000000001",	-- 464: 	lw	%r11, [%sp + 1]
"00111101011010100000000000000001",	-- 465: 	sw	%r11, [%r10 + 1]
"10000100000111010110000000000000",	-- 466: 	add	%r12, %r0, %hp
"10100111101111010000000000000011",	-- 467: 	addi	%hp, %hp, 3
"10100100000011010000101011010111",	-- 468: 	addi	%r13, %r0, read_object.2704
"00111101101011000000000000000000",	-- 469: 	sw	%r13, [%r12 + 0]
"00111101010011000000000000000010",	-- 470: 	sw	%r10, [%r12 + 2]
"00111011110010100000000000000000",	-- 471: 	lw	%r10, [%sp + 0]
"00111101010011000000000000000001",	-- 472: 	sw	%r10, [%r12 + 1]
"10000100000111010110100000000000",	-- 473: 	add	%r13, %r0, %hp
"10100111101111010000000000000010",	-- 474: 	addi	%hp, %hp, 2
"10100100000011100000101011110100",	-- 475: 	addi	%r14, %r0, read_all_object.2706
"00111101110011010000000000000000",	-- 476: 	sw	%r14, [%r13 + 0]
"00111101100011010000000000000001",	-- 477: 	sw	%r12, [%r13 + 1]
"10000100000111010110000000000000",	-- 478: 	add	%r12, %r0, %hp
"10100111101111010000000000000010",	-- 479: 	addi	%hp, %hp, 2
"10100100000011100000101100110111",	-- 480: 	addi	%r14, %r0, read_and_network.2712
"00111101110011000000000000000000",	-- 481: 	sw	%r14, [%r12 + 0]
"00111011110011100000000000000111",	-- 482: 	lw	%r14, [%sp + 7]
"00111101110011000000000000000001",	-- 483: 	sw	%r14, [%r12 + 1]
"10000100000111010111100000000000",	-- 484: 	add	%r15, %r0, %hp
"10100111101111010000000000000110",	-- 485: 	addi	%hp, %hp, 6
"10100100000100000000101101010010",	-- 486: 	addi	%r16, %r0, read_parameter.2714
"00111110000011110000000000000000",	-- 487: 	sw	%r16, [%r15 + 0]
"00111100010011110000000000000101",	-- 488: 	sw	%r2, [%r15 + 5]
"00111100111011110000000000000100",	-- 489: 	sw	%r7, [%r15 + 4]
"00111101100011110000000000000011",	-- 490: 	sw	%r12, [%r15 + 3]
"00111101101011110000000000000010",	-- 491: 	sw	%r13, [%r15 + 2]
"00111011110000100000000000001001",	-- 492: 	lw	%r2, [%sp + 9]
"00111100010011110000000000000001",	-- 493: 	sw	%r2, [%r15 + 1]
"10000100000111010011100000000000",	-- 494: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 495: 	addi	%hp, %hp, 2
"10100100000011000000101110000110",	-- 496: 	addi	%r12, %r0, solver_rect_surface.2716
"00111101100001110000000000000000",	-- 497: 	sw	%r12, [%r7 + 0]
"00111011110011000000000000001010",	-- 498: 	lw	%r12, [%sp + 10]
"00111101100001110000000000000001",	-- 499: 	sw	%r12, [%r7 + 1]
"10000100000111010110100000000000",	-- 500: 	add	%r13, %r0, %hp
"10100111101111010000000000000010",	-- 501: 	addi	%hp, %hp, 2
"10100100000100000000110000000110",	-- 502: 	addi	%r16, %r0, solver_rect.2725
"00111110000011010000000000000000",	-- 503: 	sw	%r16, [%r13 + 0]
"00111100111011010000000000000001",	-- 504: 	sw	%r7, [%r13 + 1]
"10000100000111010011100000000000",	-- 505: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 506: 	addi	%hp, %hp, 2
"10100100000100000000110001000010",	-- 507: 	addi	%r16, %r0, solver_surface.2731
"00111110000001110000000000000000",	-- 508: 	sw	%r16, [%r7 + 0]
"00111101100001110000000000000001",	-- 509: 	sw	%r12, [%r7 + 1]
"10000100000111011000000000000000",	-- 510: 	add	%r16, %r0, %hp
"10100111101111010000000000000010",	-- 511: 	addi	%hp, %hp, 2
"10100100000100010000110101011111",	-- 512: 	addi	%r17, %r0, solver_second.2750
"00111110001100000000000000000000",	-- 513: 	sw	%r17, [%r16 + 0]
"00111101100100000000000000000001",	-- 514: 	sw	%r12, [%r16 + 1]
"10000100000111011000100000000000",	-- 515: 	add	%r17, %r0, %hp
"10100111101111010000000000000101",	-- 516: 	addi	%hp, %hp, 5
"10100100000100100000110111100111",	-- 517: 	addi	%r18, %r0, solver.2756
"00111110010100010000000000000000",	-- 518: 	sw	%r18, [%r17 + 0]
"00111100111100010000000000000100",	-- 519: 	sw	%r7, [%r17 + 4]
"00111110000100010000000000000011",	-- 520: 	sw	%r16, [%r17 + 3]
"00111101101100010000000000000010",	-- 521: 	sw	%r13, [%r17 + 2]
"00111101011100010000000000000001",	-- 522: 	sw	%r11, [%r17 + 1]
"10000100000111010011100000000000",	-- 523: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 524: 	addi	%hp, %hp, 2
"10100100000011010000111000111101",	-- 525: 	addi	%r13, %r0, solver_rect_fast.2760
"00111101101001110000000000000000",	-- 526: 	sw	%r13, [%r7 + 0]
"00111101100001110000000000000001",	-- 527: 	sw	%r12, [%r7 + 1]
"10000100000111010110100000000000",	-- 528: 	add	%r13, %r0, %hp
"10100111101111010000000000000010",	-- 529: 	addi	%hp, %hp, 2
"10100100000100000000111101100011",	-- 530: 	addi	%r16, %r0, solver_surface_fast.2767
"00111110000011010000000000000000",	-- 531: 	sw	%r16, [%r13 + 0]
"00111101100011010000000000000001",	-- 532: 	sw	%r12, [%r13 + 1]
"10000100000111011000000000000000",	-- 533: 	add	%r16, %r0, %hp
"10100111101111010000000000000010",	-- 534: 	addi	%hp, %hp, 2
"10100100000100100000111110001110",	-- 535: 	addi	%r18, %r0, solver_second_fast.2773
"00111110010100000000000000000000",	-- 536: 	sw	%r18, [%r16 + 0]
"00111101100100000000000000000001",	-- 537: 	sw	%r12, [%r16 + 1]
"10000100000111011001000000000000",	-- 538: 	add	%r18, %r0, %hp
"10100111101111010000000000000101",	-- 539: 	addi	%hp, %hp, 5
"10100100000100110001000000010101",	-- 540: 	addi	%r19, %r0, solver_fast.2779
"00111110011100100000000000000000",	-- 541: 	sw	%r19, [%r18 + 0]
"00111101101100100000000000000100",	-- 542: 	sw	%r13, [%r18 + 4]
"00111110000100100000000000000011",	-- 543: 	sw	%r16, [%r18 + 3]
"00111100111100100000000000000010",	-- 544: 	sw	%r7, [%r18 + 2]
"00111101011100100000000000000001",	-- 545: 	sw	%r11, [%r18 + 1]
"10000100000111010110100000000000",	-- 546: 	add	%r13, %r0, %hp
"10100111101111010000000000000010",	-- 547: 	addi	%hp, %hp, 2
"10100100000100000001000001111111",	-- 548: 	addi	%r16, %r0, solver_surface_fast2.2783
"00111110000011010000000000000000",	-- 549: 	sw	%r16, [%r13 + 0]
"00111101100011010000000000000001",	-- 550: 	sw	%r12, [%r13 + 1]
"10000100000111011000000000000000",	-- 551: 	add	%r16, %r0, %hp
"10100111101111010000000000000010",	-- 552: 	addi	%hp, %hp, 2
"10100100000100110001000010011110",	-- 553: 	addi	%r19, %r0, solver_second_fast2.2790
"00111110011100000000000000000000",	-- 554: 	sw	%r19, [%r16 + 0]
"00111101100100000000000000000001",	-- 555: 	sw	%r12, [%r16 + 1]
"10000100000111011001100000000000",	-- 556: 	add	%r19, %r0, %hp
"10100111101111010000000000000101",	-- 557: 	addi	%hp, %hp, 5
"10100100000101000001000100010000",	-- 558: 	addi	%r20, %r0, solver_fast2.2797
"00111110100100110000000000000000",	-- 559: 	sw	%r20, [%r19 + 0]
"00111101101100110000000000000100",	-- 560: 	sw	%r13, [%r19 + 4]
"00111110000100110000000000000011",	-- 561: 	sw	%r16, [%r19 + 3]
"00111100111100110000000000000010",	-- 562: 	sw	%r7, [%r19 + 2]
"00111101011100110000000000000001",	-- 563: 	sw	%r11, [%r19 + 1]
"10000100000111010011100000000000",	-- 564: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 565: 	addi	%hp, %hp, 2
"10100100000011010001001111100001",	-- 566: 	addi	%r13, %r0, iter_setup_dirvec_constants.2809
"00111101101001110000000000000000",	-- 567: 	sw	%r13, [%r7 + 0]
"00111101011001110000000000000001",	-- 568: 	sw	%r11, [%r7 + 1]
"10000100000111010110100000000000",	-- 569: 	add	%r13, %r0, %hp
"10100111101111010000000000000011",	-- 570: 	addi	%hp, %hp, 3
"10100100000100000001010000101101",	-- 571: 	addi	%r16, %r0, setup_dirvec_constants.2812
"00111110000011010000000000000000",	-- 572: 	sw	%r16, [%r13 + 0]
"00111101010011010000000000000010",	-- 573: 	sw	%r10, [%r13 + 2]
"00111100111011010000000000000001",	-- 574: 	sw	%r7, [%r13 + 1]
"10000100000111010011100000000000",	-- 575: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 576: 	addi	%hp, %hp, 2
"10100100000100000001010000110110",	-- 577: 	addi	%r16, %r0, setup_startp_constants.2814
"00111110000001110000000000000000",	-- 578: 	sw	%r16, [%r7 + 0]
"00111101011001110000000000000001",	-- 579: 	sw	%r11, [%r7 + 1]
"10000100000111011000000000000000",	-- 580: 	add	%r16, %r0, %hp
"10100111101111010000000000000100",	-- 581: 	addi	%hp, %hp, 4
"10100100000101000001010011001111",	-- 582: 	addi	%r20, %r0, setup_startp.2817
"00111110100100000000000000000000",	-- 583: 	sw	%r20, [%r16 + 0]
"00111011110101000000000000010111",	-- 584: 	lw	%r20, [%sp + 23]
"00111110100100000000000000000011",	-- 585: 	sw	%r20, [%r16 + 3]
"00111100111100000000000000000010",	-- 586: 	sw	%r7, [%r16 + 2]
"00111101010100000000000000000001",	-- 587: 	sw	%r10, [%r16 + 1]
"10000100000111010011100000000000",	-- 588: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 589: 	addi	%hp, %hp, 2
"10100100000101010001010111010000",	-- 590: 	addi	%r21, %r0, check_all_inside.2839
"00111110101001110000000000000000",	-- 591: 	sw	%r21, [%r7 + 0]
"00111101011001110000000000000001",	-- 592: 	sw	%r11, [%r7 + 1]
"10000100000111011010100000000000",	-- 593: 	add	%r21, %r0, %hp
"10100111101111010000000000001000",	-- 594: 	addi	%hp, %hp, 8
"10100100000101100001010111110100",	-- 595: 	addi	%r22, %r0, shadow_check_and_group.2845
"00111110110101010000000000000000",	-- 596: 	sw	%r22, [%r21 + 0]
"00111110010101010000000000000111",	-- 597: 	sw	%r18, [%r21 + 7]
"00111101100101010000000000000110",	-- 598: 	sw	%r12, [%r21 + 6]
"00111101011101010000000000000101",	-- 599: 	sw	%r11, [%r21 + 5]
"00111011110101100000000000100000",	-- 600: 	lw	%r22, [%sp + 32]
"00111110110101010000000000000100",	-- 601: 	sw	%r22, [%r21 + 4]
"00111101000101010000000000000011",	-- 602: 	sw	%r8, [%r21 + 3]
"00111011110101110000000000001101",	-- 603: 	lw	%r23, [%sp + 13]
"00111110111101010000000000000010",	-- 604: 	sw	%r23, [%r21 + 2]
"00111100111101010000000000000001",	-- 605: 	sw	%r7, [%r21 + 1]
"10000100000111011100000000000000",	-- 606: 	add	%r24, %r0, %hp
"10100111101111010000000000000011",	-- 607: 	addi	%hp, %hp, 3
"10100100000110010001011001110011",	-- 608: 	addi	%r25, %r0, shadow_check_one_or_group.2848
"00111111001110000000000000000000",	-- 609: 	sw	%r25, [%r24 + 0]
"00111110101110000000000000000010",	-- 610: 	sw	%r21, [%r24 + 2]
"00111101110110000000000000000001",	-- 611: 	sw	%r14, [%r24 + 1]
"10000100000111011010100000000000",	-- 612: 	add	%r21, %r0, %hp
"10100111101111010000000000000110",	-- 613: 	addi	%hp, %hp, 6
"10100100000110010001011010010110",	-- 614: 	addi	%r25, %r0, shadow_check_one_or_matrix.2851
"00111111001101010000000000000000",	-- 615: 	sw	%r25, [%r21 + 0]
"00111110010101010000000000000101",	-- 616: 	sw	%r18, [%r21 + 5]
"00111101100101010000000000000100",	-- 617: 	sw	%r12, [%r21 + 4]
"00111111000101010000000000000011",	-- 618: 	sw	%r24, [%r21 + 3]
"00111110110101010000000000000010",	-- 619: 	sw	%r22, [%r21 + 2]
"00111110111101010000000000000001",	-- 620: 	sw	%r23, [%r21 + 1]
"10000100000111011001000000000000",	-- 621: 	add	%r18, %r0, %hp
"10100111101111010000000000001010",	-- 622: 	addi	%hp, %hp, 10
"10100100000110000001011011110111",	-- 623: 	addi	%r24, %r0, solve_each_element.2854
"00111111000100100000000000000000",	-- 624: 	sw	%r24, [%r18 + 0]
"00111011110110000000000000001100",	-- 625: 	lw	%r24, [%sp + 12]
"00111111000100100000000000001001",	-- 626: 	sw	%r24, [%r18 + 9]
"00111011110110010000000000010110",	-- 627: 	lw	%r25, [%sp + 22]
"00111111001100100000000000001000",	-- 628: 	sw	%r25, [%r18 + 8]
"00111101100100100000000000000111",	-- 629: 	sw	%r12, [%r18 + 7]
"00111110001100100000000000000110",	-- 630: 	sw	%r17, [%r18 + 6]
"00111101011100100000000000000101",	-- 631: 	sw	%r11, [%r18 + 5]
"00111011110110100000000000001011",	-- 632: 	lw	%r26, [%sp + 11]
"00111111010100100000000000000100",	-- 633: 	sw	%r26, [%r18 + 4]
"00111110111100100000000000000011",	-- 634: 	sw	%r23, [%r18 + 3]
"00111011110110110000000000001110",	-- 635: 	lw	%r27, [%sp + 14]
"00111111011100100000000000000010",	-- 636: 	sw	%r27, [%r18 + 2]
"00111100111100100000000000000001",	-- 637: 	sw	%r7, [%r18 + 1]
"10000100000111011011000000000000",	-- 638: 	add	%r22, %r0, %hp
"10100111101111010000000000000011",	-- 639: 	addi	%hp, %hp, 3
"00111101111111100000000000100011",	-- 640: 	sw	%r15, [%sp + 35]
"10100100000011110001011110100010",	-- 641: 	addi	%r15, %r0, solve_one_or_network.2858
"00111101111101100000000000000000",	-- 642: 	sw	%r15, [%r22 + 0]
"00111110010101100000000000000010",	-- 643: 	sw	%r18, [%r22 + 2]
"00111101110101100000000000000001",	-- 644: 	sw	%r14, [%r22 + 1]
"10000100000111010111100000000000",	-- 645: 	add	%r15, %r0, %hp
"10100111101111010000000000000110",	-- 646: 	addi	%hp, %hp, 6
"10100100000100100001011111000010",	-- 647: 	addi	%r18, %r0, trace_or_matrix.2862
"00111110010011110000000000000000",	-- 648: 	sw	%r18, [%r15 + 0]
"00111111000011110000000000000101",	-- 649: 	sw	%r24, [%r15 + 5]
"00111111001011110000000000000100",	-- 650: 	sw	%r25, [%r15 + 4]
"00111101100011110000000000000011",	-- 651: 	sw	%r12, [%r15 + 3]
"00111110001011110000000000000010",	-- 652: 	sw	%r17, [%r15 + 2]
"00111110110011110000000000000001",	-- 653: 	sw	%r22, [%r15 + 1]
"10000100000111011000100000000000",	-- 654: 	add	%r17, %r0, %hp
"10100111101111010000000000000100",	-- 655: 	addi	%hp, %hp, 4
"10100100000100100001100000010100",	-- 656: 	addi	%r18, %r0, judge_intersection.2866
"00111110010100010000000000000000",	-- 657: 	sw	%r18, [%r17 + 0]
"00111101111100010000000000000011",	-- 658: 	sw	%r15, [%r17 + 3]
"00111111000100010000000000000010",	-- 659: 	sw	%r24, [%r17 + 2]
"00111100010100010000000000000001",	-- 660: 	sw	%r2, [%r17 + 1]
"10000100000111010111100000000000",	-- 661: 	add	%r15, %r0, %hp
"10100111101111010000000000001010",	-- 662: 	addi	%hp, %hp, 10
"10100100000100100001100000111111",	-- 663: 	addi	%r18, %r0, solve_each_element_fast.2868
"00111110010011110000000000000000",	-- 664: 	sw	%r18, [%r15 + 0]
"00111111000011110000000000001001",	-- 665: 	sw	%r24, [%r15 + 9]
"00111110100011110000000000001000",	-- 666: 	sw	%r20, [%r15 + 8]
"00111110011011110000000000000111",	-- 667: 	sw	%r19, [%r15 + 7]
"00111101100011110000000000000110",	-- 668: 	sw	%r12, [%r15 + 6]
"00111101011011110000000000000101",	-- 669: 	sw	%r11, [%r15 + 5]
"00111111010011110000000000000100",	-- 670: 	sw	%r26, [%r15 + 4]
"00111110111011110000000000000011",	-- 671: 	sw	%r23, [%r15 + 3]
"00111111011011110000000000000010",	-- 672: 	sw	%r27, [%r15 + 2]
"00111100111011110000000000000001",	-- 673: 	sw	%r7, [%r15 + 1]
"10000100000111010011100000000000",	-- 674: 	add	%r7, %r0, %hp
"10100111101111010000000000000011",	-- 675: 	addi	%hp, %hp, 3
"10100100000100100001100011110011",	-- 676: 	addi	%r18, %r0, solve_one_or_network_fast.2872
"00111110010001110000000000000000",	-- 677: 	sw	%r18, [%r7 + 0]
"00111101111001110000000000000010",	-- 678: 	sw	%r15, [%r7 + 2]
"00111101110001110000000000000001",	-- 679: 	sw	%r14, [%r7 + 1]
"10000100000111010111000000000000",	-- 680: 	add	%r14, %r0, %hp
"10100111101111010000000000000101",	-- 681: 	addi	%hp, %hp, 5
"10100100000011110001100100010011",	-- 682: 	addi	%r15, %r0, trace_or_matrix_fast.2876
"00111101111011100000000000000000",	-- 683: 	sw	%r15, [%r14 + 0]
"00111111000011100000000000000100",	-- 684: 	sw	%r24, [%r14 + 4]
"00111110011011100000000000000011",	-- 685: 	sw	%r19, [%r14 + 3]
"00111101100011100000000000000010",	-- 686: 	sw	%r12, [%r14 + 2]
"00111100111011100000000000000001",	-- 687: 	sw	%r7, [%r14 + 1]
"10000100000111010011100000000000",	-- 688: 	add	%r7, %r0, %hp
"10100111101111010000000000000100",	-- 689: 	addi	%hp, %hp, 4
"10100100000011000001100101100011",	-- 690: 	addi	%r12, %r0, judge_intersection_fast.2880
"00111101100001110000000000000000",	-- 691: 	sw	%r12, [%r7 + 0]
"00111101110001110000000000000011",	-- 692: 	sw	%r14, [%r7 + 3]
"00111111000001110000000000000010",	-- 693: 	sw	%r24, [%r7 + 2]
"00111100010001110000000000000001",	-- 694: 	sw	%r2, [%r7 + 1]
"10000100000111010110000000000000",	-- 695: 	add	%r12, %r0, %hp
"10100111101111010000000000000011",	-- 696: 	addi	%hp, %hp, 3
"10100100000011100001100110001110",	-- 697: 	addi	%r14, %r0, get_nvector_rect.2882
"00111101110011000000000000000000",	-- 698: 	sw	%r14, [%r12 + 0]
"00111011110011100000000000001111",	-- 699: 	lw	%r14, [%sp + 15]
"00111101110011000000000000000010",	-- 700: 	sw	%r14, [%r12 + 2]
"00111111010011000000000000000001",	-- 701: 	sw	%r26, [%r12 + 1]
"10000100000111010111100000000000",	-- 702: 	add	%r15, %r0, %hp
"10100111101111010000000000000010",	-- 703: 	addi	%hp, %hp, 2
"10100100000100100001100110110100",	-- 704: 	addi	%r18, %r0, get_nvector_plane.2884
"00111110010011110000000000000000",	-- 705: 	sw	%r18, [%r15 + 0]
"00111101110011110000000000000001",	-- 706: 	sw	%r14, [%r15 + 1]
"10000100000111011001000000000000",	-- 707: 	add	%r18, %r0, %hp
"10100111101111010000000000000011",	-- 708: 	addi	%hp, %hp, 3
"10100100000100110001100111101100",	-- 709: 	addi	%r19, %r0, get_nvector_second.2886
"00111110011100100000000000000000",	-- 710: 	sw	%r19, [%r18 + 0]
"00111101110100100000000000000010",	-- 711: 	sw	%r14, [%r18 + 2]
"00111110111100100000000000000001",	-- 712: 	sw	%r23, [%r18 + 1]
"10000100000111011001100000000000",	-- 713: 	add	%r19, %r0, %hp
"10100111101111010000000000000100",	-- 714: 	addi	%hp, %hp, 4
"10100100000101000001101010110110",	-- 715: 	addi	%r20, %r0, get_nvector.2888
"00111110100100110000000000000000",	-- 716: 	sw	%r20, [%r19 + 0]
"00111110010100110000000000000011",	-- 717: 	sw	%r18, [%r19 + 3]
"00111101100100110000000000000010",	-- 718: 	sw	%r12, [%r19 + 2]
"00111101111100110000000000000001",	-- 719: 	sw	%r15, [%r19 + 1]
"10000100000111010110000000000000",	-- 720: 	add	%r12, %r0, %hp
"10100111101111010000000000000010",	-- 721: 	addi	%hp, %hp, 2
"10100100000011110001101011010011",	-- 722: 	addi	%r15, %r0, utexture.2891
"00111101111011000000000000000000",	-- 723: 	sw	%r15, [%r12 + 0]
"00111011110011110000000000010000",	-- 724: 	lw	%r15, [%sp + 16]
"00111101111011000000000000000001",	-- 725: 	sw	%r15, [%r12 + 1]
"10000100000111011001000000000000",	-- 726: 	add	%r18, %r0, %hp
"10100111101111010000000000000011",	-- 727: 	addi	%hp, %hp, 3
"10100100000101000001110011100001",	-- 728: 	addi	%r20, %r0, add_light.2894
"00111110100100100000000000000000",	-- 729: 	sw	%r20, [%r18 + 0]
"00111101111100100000000000000010",	-- 730: 	sw	%r15, [%r18 + 2]
"00111011110101000000000000010010",	-- 731: 	lw	%r20, [%sp + 18]
"00111110100100100000000000000001",	-- 732: 	sw	%r20, [%r18 + 1]
"10000100000111011011000000000000",	-- 733: 	add	%r22, %r0, %hp
"10100111101111010000000000001001",	-- 734: 	addi	%hp, %hp, 9
"00111101101111100000000000100100",	-- 735: 	sw	%r13, [%sp + 36]
"10100100000011010001110100100101",	-- 736: 	addi	%r13, %r0, trace_reflections.2898
"00111101101101100000000000000000",	-- 737: 	sw	%r13, [%r22 + 0]
"00111110101101100000000000001000",	-- 738: 	sw	%r21, [%r22 + 8]
"00111011110011010000000000100010",	-- 739: 	lw	%r13, [%sp + 34]
"00111101101101100000000000000111",	-- 740: 	sw	%r13, [%r22 + 7]
"00111100010101100000000000000110",	-- 741: 	sw	%r2, [%r22 + 6]
"00111101110101100000000000000101",	-- 742: 	sw	%r14, [%r22 + 5]
"00111100111101100000000000000100",	-- 743: 	sw	%r7, [%r22 + 4]
"00111111010101100000000000000011",	-- 744: 	sw	%r26, [%r22 + 3]
"00111111011101100000000000000010",	-- 745: 	sw	%r27, [%r22 + 2]
"00111110010101100000000000000001",	-- 746: 	sw	%r18, [%r22 + 1]
"10000100000111010110100000000000",	-- 747: 	add	%r13, %r0, %hp
"10100111101111010000000000010101",	-- 748: 	addi	%hp, %hp, 21
"10100100000010100001110110110000",	-- 749: 	addi	%r10, %r0, trace_ray.2903
"00111101010011010000000000000000",	-- 750: 	sw	%r10, [%r13 + 0]
"00111101100011010000000000010100",	-- 751: 	sw	%r12, [%r13 + 20]
"00111110110011010000000000010011",	-- 752: 	sw	%r22, [%r13 + 19]
"00111111000011010000000000010010",	-- 753: 	sw	%r24, [%r13 + 18]
"00111101111011010000000000010001",	-- 754: 	sw	%r15, [%r13 + 17]
"00111111001011010000000000010000",	-- 755: 	sw	%r25, [%r13 + 16]
"00111110101011010000000000001111",	-- 756: 	sw	%r21, [%r13 + 15]
"00111110000011010000000000001110",	-- 757: 	sw	%r16, [%r13 + 14]
"00111110100011010000000000001101",	-- 758: 	sw	%r20, [%r13 + 13]
"00111100010011010000000000001100",	-- 759: 	sw	%r2, [%r13 + 12]
"00111101011011010000000000001011",	-- 760: 	sw	%r11, [%r13 + 11]
"00111101110011010000000000001010",	-- 761: 	sw	%r14, [%r13 + 10]
"00111100001011010000000000001001",	-- 762: 	sw	%r1, [%r13 + 9]
"00111101000011010000000000001000",	-- 763: 	sw	%r8, [%r13 + 8]
"00111110001011010000000000000111",	-- 764: 	sw	%r17, [%r13 + 7]
"00111111010011010000000000000110",	-- 765: 	sw	%r26, [%r13 + 6]
"00111110111011010000000000000101",	-- 766: 	sw	%r23, [%r13 + 5]
"00111111011011010000000000000100",	-- 767: 	sw	%r27, [%r13 + 4]
"00111110011011010000000000000011",	-- 768: 	sw	%r19, [%r13 + 3]
"00111101001011010000000000000010",	-- 769: 	sw	%r9, [%r13 + 2]
"00111110010011010000000000000001",	-- 770: 	sw	%r18, [%r13 + 1]
"10000100000111010100100000000000",	-- 771: 	add	%r9, %r0, %hp
"10100111101111010000000000001101",	-- 772: 	addi	%hp, %hp, 13
"10100100000010100001111101110101",	-- 773: 	addi	%r10, %r0, trace_diffuse_ray.2909
"00111101010010010000000000000000",	-- 774: 	sw	%r10, [%r9 + 0]
"00111101100010010000000000001100",	-- 775: 	sw	%r12, [%r9 + 12]
"00111101111010010000000000001011",	-- 776: 	sw	%r15, [%r9 + 11]
"00111110101010010000000000001010",	-- 777: 	sw	%r21, [%r9 + 10]
"00111100010010010000000000001001",	-- 778: 	sw	%r2, [%r9 + 9]
"00111101011010010000000000001000",	-- 779: 	sw	%r11, [%r9 + 8]
"00111101110010010000000000000111",	-- 780: 	sw	%r14, [%r9 + 7]
"00111101000010010000000000000110",	-- 781: 	sw	%r8, [%r9 + 6]
"00111100111010010000000000000101",	-- 782: 	sw	%r7, [%r9 + 5]
"00111110111010010000000000000100",	-- 783: 	sw	%r23, [%r9 + 4]
"00111111011010010000000000000011",	-- 784: 	sw	%r27, [%r9 + 3]
"00111110011010010000000000000010",	-- 785: 	sw	%r19, [%r9 + 2]
"00111011110000100000000000010001",	-- 786: 	lw	%r2, [%sp + 17]
"00111100010010010000000000000001",	-- 787: 	sw	%r2, [%r9 + 1]
"10000100000111010011100000000000",	-- 788: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 789: 	addi	%hp, %hp, 2
"10100100000010100001111111101110",	-- 790: 	addi	%r10, %r0, iter_trace_diffuse_rays.2912
"00111101010001110000000000000000",	-- 791: 	sw	%r10, [%r7 + 0]
"00111101001001110000000000000001",	-- 792: 	sw	%r9, [%r7 + 1]
"10000100000111010100100000000000",	-- 793: 	add	%r9, %r0, %hp
"10100111101111010000000000000011",	-- 794: 	addi	%hp, %hp, 3
"10100100000010100010000000111001",	-- 795: 	addi	%r10, %r0, trace_diffuse_rays.2917
"00111101010010010000000000000000",	-- 796: 	sw	%r10, [%r9 + 0]
"00111110000010010000000000000010",	-- 797: 	sw	%r16, [%r9 + 2]
"00111100111010010000000000000001",	-- 798: 	sw	%r7, [%r9 + 1]
"10000100000111010011100000000000",	-- 799: 	add	%r7, %r0, %hp
"10100111101111010000000000000011",	-- 800: 	addi	%hp, %hp, 3
"10100100000010100010000001001110",	-- 801: 	addi	%r10, %r0, trace_diffuse_ray_80percent.2921
"00111101010001110000000000000000",	-- 802: 	sw	%r10, [%r7 + 0]
"00111101001001110000000000000010",	-- 803: 	sw	%r9, [%r7 + 2]
"00111011110010100000000000011101",	-- 804: 	lw	%r10, [%sp + 29]
"00111101010001110000000000000001",	-- 805: 	sw	%r10, [%r7 + 1]
"10000100000111010110000000000000",	-- 806: 	add	%r12, %r0, %hp
"10100111101111010000000000000100",	-- 807: 	addi	%hp, %hp, 4
"10100100000011100010000010101001",	-- 808: 	addi	%r14, %r0, calc_diffuse_using_1point.2925
"00111101110011000000000000000000",	-- 809: 	sw	%r14, [%r12 + 0]
"00111100111011000000000000000011",	-- 810: 	sw	%r7, [%r12 + 3]
"00111110100011000000000000000010",	-- 811: 	sw	%r20, [%r12 + 2]
"00111100010011000000000000000001",	-- 812: 	sw	%r2, [%r12 + 1]
"10000100000111010011100000000000",	-- 813: 	add	%r7, %r0, %hp
"10100111101111010000000000000011",	-- 814: 	addi	%hp, %hp, 3
"10100100000011100010000011111000",	-- 815: 	addi	%r14, %r0, calc_diffuse_using_5points.2928
"00111101110001110000000000000000",	-- 816: 	sw	%r14, [%r7 + 0]
"00111110100001110000000000000010",	-- 817: 	sw	%r20, [%r7 + 2]
"00111100010001110000000000000001",	-- 818: 	sw	%r2, [%r7 + 1]
"10000100000111010111000000000000",	-- 819: 	add	%r14, %r0, %hp
"10100111101111010000000000000010",	-- 820: 	addi	%hp, %hp, 2
"10100100000011110010000110000000",	-- 821: 	addi	%r15, %r0, do_without_neighbors.2934
"00111101111011100000000000000000",	-- 822: 	sw	%r15, [%r14 + 0]
"00111101100011100000000000000001",	-- 823: 	sw	%r12, [%r14 + 1]
"10000100000111010110000000000000",	-- 824: 	add	%r12, %r0, %hp
"10100111101111010000000000000010",	-- 825: 	addi	%hp, %hp, 2
"10100100000011110010000110101110",	-- 826: 	addi	%r15, %r0, neighbors_exist.2937
"00111101111011000000000000000000",	-- 827: 	sw	%r15, [%r12 + 0]
"00111011110011110000000000010011",	-- 828: 	lw	%r15, [%sp + 19]
"00111101111011000000000000000001",	-- 829: 	sw	%r15, [%r12 + 1]
"10000100000111011000000000000000",	-- 830: 	add	%r16, %r0, %hp
"10100111101111010000000000000011",	-- 831: 	addi	%hp, %hp, 3
"10100100000100010010001000100110",	-- 832: 	addi	%r17, %r0, try_exploit_neighbors.2950
"00111110001100000000000000000000",	-- 833: 	sw	%r17, [%r16 + 0]
"00111101110100000000000000000010",	-- 834: 	sw	%r14, [%r16 + 2]
"00111100111100000000000000000001",	-- 835: 	sw	%r7, [%r16 + 1]
"10000100000111010011100000000000",	-- 836: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 837: 	addi	%hp, %hp, 2
"10100100000100010010001001111001",	-- 838: 	addi	%r17, %r0, write_ppm_header.2957
"00111110001001110000000000000000",	-- 839: 	sw	%r17, [%r7 + 0]
"00111101111001110000000000000001",	-- 840: 	sw	%r15, [%r7 + 1]
"10000100000111011000100000000000",	-- 841: 	add	%r17, %r0, %hp
"10100111101111010000000000000010",	-- 842: 	addi	%hp, %hp, 2
"10100100000100100010001011000010",	-- 843: 	addi	%r18, %r0, write_rgb.2961
"00111110010100010000000000000000",	-- 844: 	sw	%r18, [%r17 + 0]
"00111110100100010000000000000001",	-- 845: 	sw	%r20, [%r17 + 1]
"10000100000111011001000000000000",	-- 846: 	add	%r18, %r0, %hp
"10100111101111010000000000000100",	-- 847: 	addi	%hp, %hp, 4
"10100100000100110010001011101100",	-- 848: 	addi	%r19, %r0, pretrace_diffuse_rays.2963
"00111110011100100000000000000000",	-- 849: 	sw	%r19, [%r18 + 0]
"00111101001100100000000000000011",	-- 850: 	sw	%r9, [%r18 + 3]
"00111101010100100000000000000010",	-- 851: 	sw	%r10, [%r18 + 2]
"00111100010100100000000000000001",	-- 852: 	sw	%r2, [%r18 + 1]
"10000100000111010001000000000000",	-- 853: 	add	%r2, %r0, %hp
"10100111101111010000000000001010",	-- 854: 	addi	%hp, %hp, 10
"10100100000010010010001101010011",	-- 855: 	addi	%r9, %r0, pretrace_pixels.2966
"00111101001000100000000000000000",	-- 856: 	sw	%r9, [%r2 + 0]
"00111100011000100000000000001001",	-- 857: 	sw	%r3, [%r2 + 9]
"00111101101000100000000000001000",	-- 858: 	sw	%r13, [%r2 + 8]
"00111111001000100000000000000111",	-- 859: 	sw	%r25, [%r2 + 7]
"00111100110000100000000000000110",	-- 860: 	sw	%r6, [%r2 + 6]
"00111011110000110000000000010101",	-- 861: 	lw	%r3, [%sp + 21]
"00111100011000100000000000000101",	-- 862: 	sw	%r3, [%r2 + 5]
"00111110100000100000000000000100",	-- 863: 	sw	%r20, [%r2 + 4]
"00111011110001100000000000011011",	-- 864: 	lw	%r6, [%sp + 27]
"00111100110000100000000000000011",	-- 865: 	sw	%r6, [%r2 + 3]
"00111110010000100000000000000010",	-- 866: 	sw	%r18, [%r2 + 2]
"00111011110001100000000000010100",	-- 867: 	lw	%r6, [%sp + 20]
"00111100110000100000000000000001",	-- 868: 	sw	%r6, [%r2 + 1]
"10000100000111010100100000000000",	-- 869: 	add	%r9, %r0, %hp
"10100111101111010000000000000111",	-- 870: 	addi	%hp, %hp, 7
"10100100000011010010010000000010",	-- 871: 	addi	%r13, %r0, pretrace_line.2973
"00111101101010010000000000000000",	-- 872: 	sw	%r13, [%r9 + 0]
"00111100100010010000000000000110",	-- 873: 	sw	%r4, [%r9 + 6]
"00111100101010010000000000000101",	-- 874: 	sw	%r5, [%r9 + 5]
"00111100011010010000000000000100",	-- 875: 	sw	%r3, [%r9 + 4]
"00111100010010010000000000000011",	-- 876: 	sw	%r2, [%r9 + 3]
"00111101111010010000000000000010",	-- 877: 	sw	%r15, [%r9 + 2]
"00111100110010010000000000000001",	-- 878: 	sw	%r6, [%r9 + 1]
"10000100000111010001000000000000",	-- 879: 	add	%r2, %r0, %hp
"10100111101111010000000000000111",	-- 880: 	addi	%hp, %hp, 7
"10100100000001000010010001000111",	-- 881: 	addi	%r4, %r0, scan_pixel.2977
"00111100100000100000000000000000",	-- 882: 	sw	%r4, [%r2 + 0]
"00111110001000100000000000000110",	-- 883: 	sw	%r17, [%r2 + 6]
"00111110000000100000000000000101",	-- 884: 	sw	%r16, [%r2 + 5]
"00111110100000100000000000000100",	-- 885: 	sw	%r20, [%r2 + 4]
"00111101100000100000000000000011",	-- 886: 	sw	%r12, [%r2 + 3]
"00111101111000100000000000000010",	-- 887: 	sw	%r15, [%r2 + 2]
"00111101110000100000000000000001",	-- 888: 	sw	%r14, [%r2 + 1]
"10000100000111010010000000000000",	-- 889: 	add	%r4, %r0, %hp
"10100111101111010000000000000100",	-- 890: 	addi	%hp, %hp, 4
"10100100000001010010010010100101",	-- 891: 	addi	%r5, %r0, scan_line.2983
"00111100101001000000000000000000",	-- 892: 	sw	%r5, [%r4 + 0]
"00111100010001000000000000000011",	-- 893: 	sw	%r2, [%r4 + 3]
"00111101001001000000000000000010",	-- 894: 	sw	%r9, [%r4 + 2]
"00111101111001000000000000000001",	-- 895: 	sw	%r15, [%r4 + 1]
"10000100000111010001000000000000",	-- 896: 	add	%r2, %r0, %hp
"10100111101111010000000000000010",	-- 897: 	addi	%hp, %hp, 2
"10100100000001010010010110011000",	-- 898: 	addi	%r5, %r0, create_pixelline.2996
"00111100101000100000000000000000",	-- 899: 	sw	%r5, [%r2 + 0]
"00111101111000100000000000000001",	-- 900: 	sw	%r15, [%r2 + 1]
"10000100000111010010100000000000",	-- 901: 	add	%r5, %r0, %hp
"10100111101111010000000000000010",	-- 902: 	addi	%hp, %hp, 2
"10100100000011000010010111100000",	-- 903: 	addi	%r12, %r0, calc_dirvec.3003
"00111101100001010000000000000000",	-- 904: 	sw	%r12, [%r5 + 0]
"00111101010001010000000000000001",	-- 905: 	sw	%r10, [%r5 + 1]
"10000100000111010110000000000000",	-- 906: 	add	%r12, %r0, %hp
"10100111101111010000000000000010",	-- 907: 	addi	%hp, %hp, 2
"10100100000011010010011011100011",	-- 908: 	addi	%r13, %r0, calc_dirvecs.3011
"00111101101011000000000000000000",	-- 909: 	sw	%r13, [%r12 + 0]
"00111100101011000000000000000001",	-- 910: 	sw	%r5, [%r12 + 1]
"10000100000111010010100000000000",	-- 911: 	add	%r5, %r0, %hp
"10100111101111010000000000000010",	-- 912: 	addi	%hp, %hp, 2
"10100100000011010010011100111001",	-- 913: 	addi	%r13, %r0, calc_dirvec_rows.3016
"00111101101001010000000000000000",	-- 914: 	sw	%r13, [%r5 + 0]
"00111101100001010000000000000001",	-- 915: 	sw	%r12, [%r5 + 1]
"10000100000111010110000000000000",	-- 916: 	add	%r12, %r0, %hp
"10100111101111010000000000000010",	-- 917: 	addi	%hp, %hp, 2
"10100100000011010010011101101011",	-- 918: 	addi	%r13, %r0, create_dirvec.3020
"00111101101011000000000000000000",	-- 919: 	sw	%r13, [%r12 + 0]
"00111011110011010000000000000000",	-- 920: 	lw	%r13, [%sp + 0]
"00111101101011000000000000000001",	-- 921: 	sw	%r13, [%r12 + 1]
"10000100000111010111000000000000",	-- 922: 	add	%r14, %r0, %hp
"10100111101111010000000000000010",	-- 923: 	addi	%hp, %hp, 2
"10100100000100000010011110001000",	-- 924: 	addi	%r16, %r0, create_dirvec_elements.3022
"00111110000011100000000000000000",	-- 925: 	sw	%r16, [%r14 + 0]
"00111101100011100000000000000001",	-- 926: 	sw	%r12, [%r14 + 1]
"10000100000111011000000000000000",	-- 927: 	add	%r16, %r0, %hp
"10100111101111010000000000000100",	-- 928: 	addi	%hp, %hp, 4
"10100100000100010010011110100000",	-- 929: 	addi	%r17, %r0, create_dirvecs.3025
"00111110001100000000000000000000",	-- 930: 	sw	%r17, [%r16 + 0]
"00111101010100000000000000000011",	-- 931: 	sw	%r10, [%r16 + 3]
"00111101110100000000000000000010",	-- 932: 	sw	%r14, [%r16 + 2]
"00111101100100000000000000000001",	-- 933: 	sw	%r12, [%r16 + 1]
"10000100000111010111000000000000",	-- 934: 	add	%r14, %r0, %hp
"10100111101111010000000000000010",	-- 935: 	addi	%hp, %hp, 2
"10100100000100010010011111001111",	-- 936: 	addi	%r17, %r0, init_dirvec_constants.3027
"00111110001011100000000000000000",	-- 937: 	sw	%r17, [%r14 + 0]
"00111011110100010000000000100100",	-- 938: 	lw	%r17, [%sp + 36]
"00111110001011100000000000000001",	-- 939: 	sw	%r17, [%r14 + 1]
"10000100000111011001000000000000",	-- 940: 	add	%r18, %r0, %hp
"10100111101111010000000000000011",	-- 941: 	addi	%hp, %hp, 3
"10100100000100110010011111100111",	-- 942: 	addi	%r19, %r0, init_vecset_constants.3030
"00111110011100100000000000000000",	-- 943: 	sw	%r19, [%r18 + 0]
"00111101110100100000000000000010",	-- 944: 	sw	%r14, [%r18 + 2]
"00111101010100100000000000000001",	-- 945: 	sw	%r10, [%r18 + 1]
"10000100000111010101000000000000",	-- 946: 	add	%r10, %r0, %hp
"10100111101111010000000000000100",	-- 947: 	addi	%hp, %hp, 4
"10100100000011100010100000000000",	-- 948: 	addi	%r14, %r0, init_dirvecs.3032
"00111101110010100000000000000000",	-- 949: 	sw	%r14, [%r10 + 0]
"00111110010010100000000000000011",	-- 950: 	sw	%r18, [%r10 + 3]
"00111110000010100000000000000010",	-- 951: 	sw	%r16, [%r10 + 2]
"00111100101010100000000000000001",	-- 952: 	sw	%r5, [%r10 + 1]
"10000100000111010010100000000000",	-- 953: 	add	%r5, %r0, %hp
"10100111101111010000000000000100",	-- 954: 	addi	%hp, %hp, 4
"10100100000011100010100000011100",	-- 955: 	addi	%r14, %r0, add_reflection.3034
"00111101110001010000000000000000",	-- 956: 	sw	%r14, [%r5 + 0]
"00111110001001010000000000000011",	-- 957: 	sw	%r17, [%r5 + 3]
"00111011110011100000000000100010",	-- 958: 	lw	%r14, [%sp + 34]
"00111101110001010000000000000010",	-- 959: 	sw	%r14, [%r5 + 2]
"00111101100001010000000000000001",	-- 960: 	sw	%r12, [%r5 + 1]
"10000100000111010110000000000000",	-- 961: 	add	%r12, %r0, %hp
"10100111101111010000000000000100",	-- 962: 	addi	%hp, %hp, 4
"10100100000011100010100001010000",	-- 963: 	addi	%r14, %r0, setup_rect_reflection.3041
"00111101110011000000000000000000",	-- 964: 	sw	%r14, [%r12 + 0]
"00111100001011000000000000000011",	-- 965: 	sw	%r1, [%r12 + 3]
"00111101000011000000000000000010",	-- 966: 	sw	%r8, [%r12 + 2]
"00111100101011000000000000000001",	-- 967: 	sw	%r5, [%r12 + 1]
"10000100000111010111000000000000",	-- 968: 	add	%r14, %r0, %hp
"10100111101111010000000000000100",	-- 969: 	addi	%hp, %hp, 4
"10100100000100000010100011010000",	-- 970: 	addi	%r16, %r0, setup_surface_reflection.3044
"00111110000011100000000000000000",	-- 971: 	sw	%r16, [%r14 + 0]
"00111100001011100000000000000011",	-- 972: 	sw	%r1, [%r14 + 3]
"00111101000011100000000000000010",	-- 973: 	sw	%r8, [%r14 + 2]
"00111100101011100000000000000001",	-- 974: 	sw	%r5, [%r14 + 1]
"10000100000111010000100000000000",	-- 975: 	add	%r1, %r0, %hp
"10100111101111010000000000000100",	-- 976: 	addi	%hp, %hp, 4
"10100100000001010010100101000110",	-- 977: 	addi	%r5, %r0, setup_reflections.3047
"00111100101000010000000000000000",	-- 978: 	sw	%r5, [%r1 + 0]
"00111101110000010000000000000011",	-- 979: 	sw	%r14, [%r1 + 3]
"00111101100000010000000000000010",	-- 980: 	sw	%r12, [%r1 + 2]
"00111101011000010000000000000001",	-- 981: 	sw	%r11, [%r1 + 1]
"10000100000111011101100000000000",	-- 982: 	add	%r27, %r0, %hp
"10100111101111010000000000001111",	-- 983: 	addi	%hp, %hp, 15
"10100100000001010010100110000000",	-- 984: 	addi	%r5, %r0, rt.3049
"00111100101110110000000000000000",	-- 985: 	sw	%r5, [%r27 + 0]
"00111100111110110000000000001110",	-- 986: 	sw	%r7, [%r27 + 14]
"00111100001110110000000000001101",	-- 987: 	sw	%r1, [%r27 + 13]
"00111110001110110000000000001100",	-- 988: 	sw	%r17, [%r27 + 12]
"00111100011110110000000000001011",	-- 989: 	sw	%r3, [%r27 + 11]
"00111100100110110000000000001010",	-- 990: 	sw	%r4, [%r27 + 10]
"00111011110000010000000000100011",	-- 991: 	lw	%r1, [%sp + 35]
"00111100001110110000000000001001",	-- 992: 	sw	%r1, [%r27 + 9]
"00111101001110110000000000001000",	-- 993: 	sw	%r9, [%r27 + 8]
"00111101101110110000000000000111",	-- 994: 	sw	%r13, [%r27 + 7]
"00111011110000010000000000100000",	-- 995: 	lw	%r1, [%sp + 32]
"00111100001110110000000000000110",	-- 996: 	sw	%r1, [%r27 + 6]
"00111101000110110000000000000101",	-- 997: 	sw	%r8, [%r27 + 5]
"00111101010110110000000000000100",	-- 998: 	sw	%r10, [%r27 + 4]
"00111101111110110000000000000011",	-- 999: 	sw	%r15, [%r27 + 3]
"00111100110110110000000000000010",	-- 1000: 	sw	%r6, [%r27 + 2]
"00111100010110110000000000000001",	-- 1001: 	sw	%r2, [%r27 + 1]
"11001100000000010000000010000000",	-- 1002: 	lli	%r1, 128
"11001100000000100000000010000000",	-- 1003: 	lli	%r2, 128
"00111111111111100000000000100101",	-- 1004: 	sw	%ra, [%sp + 37]
"00111011011110100000000000000000",	-- 1005: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100110",	-- 1006: 	addi	%sp, %sp, 38
"01010011010000000000000000000000",	-- 1007: 	jalr	%r26
"10101011110111100000000000100110",	-- 1008: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 1009: 	lw	%ra, [%sp + 37]
"11001100000000010000000000000000",	-- 1010: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 1011: 	jr	%ra
	-- halt:
"11111100000000000000000000000000",	-- 1012: 	halt
	-- div10_sub.6209:
"11001100000000110000000000001010",	-- 1013: 	lli	%r3, 10
"00110000011000010000000000000110",	-- 1014: 	bgt	%r3, %r1, bgt_else.8923
"11001100000000110000000000001010",	-- 1015: 	lli	%r3, 10
"10001000001000110000100000000000",	-- 1016: 	sub	%r1, %r1, %r3
"11001100000000110000000000000001",	-- 1017: 	lli	%r3, 1
"10000100010000110001000000000000",	-- 1018: 	add	%r2, %r2, %r3
"01010100000000000000001111110101",	-- 1019: 	j	div10_sub.6209
	-- bgt_else.8923:
"10000100000000100000100000000000",	-- 1020: 	add	%r1, %r0, %r2
"01001111111000000000000000000000",	-- 1021: 	jr	%ra
	-- div10.6193:
"11001100000000100000000000000000",	-- 1022: 	lli	%r2, 0
"01010100000000000000001111110101",	-- 1023: 	j	div10_sub.6209
	-- print_int.2514:
"11001100000000100000000000000000",	-- 1024: 	lli	%r2, 0
"00110000010000010000000000011010",	-- 1025: 	bgt	%r2, %r1, bgt_else.8924
"11001100000000100000000000001010",	-- 1026: 	lli	%r2, 10
"00110000010000010000000000010101",	-- 1027: 	bgt	%r2, %r1, bgt_else.8925
"00111100001111100000000000000000",	-- 1028: 	sw	%r1, [%sp + 0]
"00111111111111100000000000000001",	-- 1029: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 1030: 	addi	%sp, %sp, 2
"01011000000000000000001111111110",	-- 1031: 	jal	div10.6193
"10101011110111100000000000000010",	-- 1032: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 1033: 	lw	%ra, [%sp + 1]
"00111100001111100000000000000001",	-- 1034: 	sw	%r1, [%sp + 1]
"00111111111111100000000000000010",	-- 1035: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1036: 	addi	%sp, %sp, 3
"01011000000000000000010000000000",	-- 1037: 	jal	print_int.2514
"10101011110111100000000000000011",	-- 1038: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1039: 	lw	%ra, [%sp + 2]
"11001100000000010000000000001010",	-- 1040: 	lli	%r1, 10
"00111011110000100000000000000001",	-- 1041: 	lw	%r2, [%sp + 1]
"10001100010000010000100000000000",	-- 1042: 	mul	%r1, %r2, %r1
"00111011110000100000000000000000",	-- 1043: 	lw	%r2, [%sp + 0]
"10001000010000010000100000000000",	-- 1044: 	sub	%r1, %r2, %r1
"11001100000000100000000000110000",	-- 1045: 	lli	%r2, 48
"10000100001000100000100000000000",	-- 1046: 	add	%r1, %r1, %r2
"01010100000000000010101000011000",	-- 1047: 	j	yj_print_char
	-- bgt_else.8925:
"11001100000000100000000000110000",	-- 1048: 	lli	%r2, 48
"10000100001000100000100000000000",	-- 1049: 	add	%r1, %r1, %r2
"01010100000000000010101000011000",	-- 1050: 	j	yj_print_char
	-- bgt_else.8924:
"11001100000000100000000000101101",	-- 1051: 	lli	%r2, 45
"00111100001111100000000000000000",	-- 1052: 	sw	%r1, [%sp + 0]
"10000100000000100000100000000000",	-- 1053: 	add	%r1, %r0, %r2
"00111111111111100000000000000010",	-- 1054: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1055: 	addi	%sp, %sp, 3
"01011000000000000010101000011000",	-- 1056: 	jal	yj_print_char
"10101011110111100000000000000011",	-- 1057: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1058: 	lw	%ra, [%sp + 2]
"00111011110000010000000000000000",	-- 1059: 	lw	%r1, [%sp + 0]
"10001000000000010000100000000000",	-- 1060: 	sub	%r1, %r0, %r1
"01010100000000000000010000000000",	-- 1061: 	j	print_int.2514
	-- calc_sin.6160:
"00010100000000011010101011000001",	-- 1062: 	llif	%f1, -0.166667
"00010000000000011011111000101010",	-- 1063: 	lhif	%f1, -0.166667
"00010100000000101000011100100011",	-- 1064: 	llif	%f2, 0.008333
"00010000000000100011110000001000",	-- 1065: 	lhif	%f2, 0.008333
"00010100000000111001111000111000",	-- 1066: 	llif	%f3, -0.000198
"00010000000000111011100101001111",	-- 1067: 	lhif	%f3, -0.000198
"00010100000001000101001110011100",	-- 1068: 	llif	%f4, 0.000003
"00010000000001000011011001001001",	-- 1069: 	lhif	%f4, 0.000003
"00010100000001010000000000000000",	-- 1070: 	llif	%f5, 0.000000
"00010000000001010000000000000000",	-- 1071: 	lhif	%f5, 0.000000
"00010100000001100000000000000000",	-- 1072: 	llif	%f6, 0.000000
"00010000000001100000000000000000",	-- 1073: 	lhif	%f6, 0.000000
"11101000000000000011100000000000",	-- 1074: 	mulf	%f7, %f0, %f0
"11101000111000000100000000000000",	-- 1075: 	mulf	%f8, %f7, %f0
"11101000111001100011000000000000",	-- 1076: 	mulf	%f6, %f7, %f6
"11100000101001100010100000000000",	-- 1077: 	addf	%f5, %f5, %f6
"11101000111001010010100000000000",	-- 1078: 	mulf	%f5, %f7, %f5
"11100000100001010010000000000000",	-- 1079: 	addf	%f4, %f4, %f5
"11101000111001000010000000000000",	-- 1080: 	mulf	%f4, %f7, %f4
"11100000011001000001100000000000",	-- 1081: 	addf	%f3, %f3, %f4
"11101000111000110001100000000000",	-- 1082: 	mulf	%f3, %f7, %f3
"11100000010000110001000000000000",	-- 1083: 	addf	%f2, %f2, %f3
"11101000111000100001000000000000",	-- 1084: 	mulf	%f2, %f7, %f2
"11100000001000100000100000000000",	-- 1085: 	addf	%f1, %f1, %f2
"11101001000000010000100000000000",	-- 1086: 	mulf	%f1, %f8, %f1
"11100000000000010000000000000000",	-- 1087: 	addf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 1088: 	jr	%ra
	-- sinf__.6162:
"00010100000000010000111111011000",	-- 1089: 	llif	%f1, 1.570796
"00010000000000010011111111001001",	-- 1090: 	lhif	%f1, 1.570796
"00010100000000100000111111011100",	-- 1091: 	llif	%f2, 3.141593
"00010000000000100100000001001001",	-- 1092: 	lhif	%f2, 3.141593
"00010100000000110000111111011010",	-- 1093: 	llif	%f3, 6.283185
"00010000000000110100000011001001",	-- 1094: 	lhif	%f3, 6.283185
"00100000000000110000000000001110",	-- 1095: 	bgtf	%f0, %f3, bgtf_else.8926
"00100000000000100000000000000101",	-- 1096: 	bgtf	%f0, %f2, bgtf_else.8927
"00100000000000010000000000000010",	-- 1097: 	bgtf	%f0, %f1, bgtf_else.8928
"01010100000000000000010000100110",	-- 1098: 	j	calc_sin.6160
	-- bgtf_else.8928:
"11100100010000000000000000000000",	-- 1099: 	subf	%f0, %f2, %f0
"01010100000000000000010001000001",	-- 1100: 	j	sinf__.6162
	-- bgtf_else.8927:
"11100100000000100000000000000000",	-- 1101: 	subf	%f0, %f0, %f2
"00111111111111100000000000000000",	-- 1102: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 1103: 	addi	%sp, %sp, 1
"01011000000000000000010001000001",	-- 1104: 	jal	sinf__.6162
"10101011110111100000000000000001",	-- 1105: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 1106: 	lw	%ra, [%sp + 0]
"00011000000000000000000000000000",	-- 1107: 	negf	%f0, %f0
"01001111111000000000000000000000",	-- 1108: 	jr	%ra
	-- bgtf_else.8926:
"11100100000000110000000000000000",	-- 1109: 	subf	%f0, %f0, %f3
"01010100000000000000010001000001",	-- 1110: 	j	sinf__.6162
	-- sin.2516:
"00010100000000010000000000000000",	-- 1111: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 1112: 	lhif	%f1, 0.000000
"00100000001000000000000000000010",	-- 1113: 	bgtf	%f1, %f0, bgtf_else.8929
"01010100000000000000010001000001",	-- 1114: 	j	sinf__.6162
	-- bgtf_else.8929:
"00011000000000000000000000000000",	-- 1115: 	negf	%f0, %f0
"00111111111111100000000000000000",	-- 1116: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 1117: 	addi	%sp, %sp, 1
"01011000000000000000010001000001",	-- 1118: 	jal	sinf__.6162
"10101011110111100000000000000001",	-- 1119: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 1120: 	lw	%ra, [%sp + 0]
"00011000000000000000000000000000",	-- 1121: 	negf	%f0, %f0
"01001111111000000000000000000000",	-- 1122: 	jr	%ra
	-- calc_cos.6127:
"00010100000000011010101100000100",	-- 1123: 	llif	%f1, 0.041667
"00010000000000010011110100101010",	-- 1124: 	lhif	%f1, 0.041667
"00010100000000100000111100011011",	-- 1125: 	llif	%f2, -0.001389
"00010000000000101011101010110110",	-- 1126: 	lhif	%f2, -0.001389
"00010100000000111011011100010111",	-- 1127: 	llif	%f3, 0.000025
"00010000000000110011011111010001",	-- 1128: 	lhif	%f3, 0.000025
"00010100000001000000000000000000",	-- 1129: 	llif	%f4, -0.000000
"00010000000001001000000000000000",	-- 1130: 	lhif	%f4, -0.000000
"00010100000001010000000000000000",	-- 1131: 	llif	%f5, -0.000000
"00010000000001011000000000000000",	-- 1132: 	lhif	%f5, -0.000000
"11101000000000000000000000000000",	-- 1133: 	mulf	%f0, %f0, %f0
"11101000000001010010100000000000",	-- 1134: 	mulf	%f5, %f0, %f5
"11100000100001010010000000000000",	-- 1135: 	addf	%f4, %f4, %f5
"11101000000001000010000000000000",	-- 1136: 	mulf	%f4, %f0, %f4
"11100000011001000001100000000000",	-- 1137: 	addf	%f3, %f3, %f4
"11101000000000110001100000000000",	-- 1138: 	mulf	%f3, %f0, %f3
"11100000010000110001000000000000",	-- 1139: 	addf	%f2, %f2, %f3
"11101000000000100001000000000000",	-- 1140: 	mulf	%f2, %f0, %f2
"11100000001000100000100000000000",	-- 1141: 	addf	%f1, %f1, %f2
"11101000000000010000100000000000",	-- 1142: 	mulf	%f1, %f0, %f1
"00010100000000100000000000000000",	-- 1143: 	llif	%f2, 1.000000
"00010000000000100011111110000000",	-- 1144: 	lhif	%f2, 1.000000
"00010100000000110000000000000000",	-- 1145: 	llif	%f3, 0.500000
"00010000000000110011111100000000",	-- 1146: 	lhif	%f3, 0.500000
"11101000011000000001100000000000",	-- 1147: 	mulf	%f3, %f3, %f0
"11100100010000110001000000000000",	-- 1148: 	subf	%f2, %f2, %f3
"11101000000000010000000000000000",	-- 1149: 	mulf	%f0, %f0, %f1
"11100000010000000000000000000000",	-- 1150: 	addf	%f0, %f2, %f0
"01001111111000000000000000000000",	-- 1151: 	jr	%ra
	-- cosf__.6129:
"00010100000000010000111111011000",	-- 1152: 	llif	%f1, 1.570796
"00010000000000010011111111001001",	-- 1153: 	lhif	%f1, 1.570796
"00010100000000100000111111011100",	-- 1154: 	llif	%f2, 3.141593
"00010000000000100100000001001001",	-- 1155: 	lhif	%f2, 3.141593
"00010100000000110000111111011010",	-- 1156: 	llif	%f3, 6.283185
"00010000000000110100000011001001",	-- 1157: 	lhif	%f3, 6.283185
"00100000000000110000000000001110",	-- 1158: 	bgtf	%f0, %f3, bgtf_else.8930
"00100000000000100000000000000101",	-- 1159: 	bgtf	%f0, %f2, bgtf_else.8931
"00100000000000010000000000000010",	-- 1160: 	bgtf	%f0, %f1, bgtf_else.8932
"01010100000000000000010001100011",	-- 1161: 	j	calc_cos.6127
	-- bgtf_else.8932:
"11100100010000000000000000000000",	-- 1162: 	subf	%f0, %f2, %f0
"01010100000000000000010010000000",	-- 1163: 	j	cosf__.6129
	-- bgtf_else.8931:
"11100100000000100000000000000000",	-- 1164: 	subf	%f0, %f0, %f2
"00111111111111100000000000000000",	-- 1165: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 1166: 	addi	%sp, %sp, 1
"01011000000000000000010010000000",	-- 1167: 	jal	cosf__.6129
"10101011110111100000000000000001",	-- 1168: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 1169: 	lw	%ra, [%sp + 0]
"00011000000000000000000000000000",	-- 1170: 	negf	%f0, %f0
"01001111111000000000000000000000",	-- 1171: 	jr	%ra
	-- bgtf_else.8930:
"11100100000000110000000000000000",	-- 1172: 	subf	%f0, %f0, %f3
"01010100000000000000010010000000",	-- 1173: 	j	cosf__.6129
	-- cos.2518:
"00010100000000010000000000000000",	-- 1174: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 1175: 	lhif	%f1, 0.000000
"00100000001000000000000000000010",	-- 1176: 	bgtf	%f1, %f0, bgtf_else.8933
"01010100000000000000010010000000",	-- 1177: 	j	cosf__.6129
	-- bgtf_else.8933:
"00011000000000000000000000000000",	-- 1178: 	negf	%f0, %f0
"01010100000000000000010010000000",	-- 1179: 	j	cosf__.6129
	-- atan.2520:
"10110000000111100000000000000000",	-- 1180: 	sf	%f0, [%sp + 0]
"00111111111111100000000000000001",	-- 1181: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 1182: 	addi	%sp, %sp, 2
"01011000000000000010101001001101",	-- 1183: 	jal	yj_fabs
"10101011110111100000000000000010",	-- 1184: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 1185: 	lw	%ra, [%sp + 1]
"00010100000000011001100110011010",	-- 1186: 	llif	%f1, 0.150000
"00010000000000010011111000011001",	-- 1187: 	lhif	%f1, 0.150000
"00100000000000010000000000010011",	-- 1188: 	bgtf	%f0, %f1, bgtf_else.8934
"10010011110000000000000000000000",	-- 1189: 	lf	%f0, [%sp + 0]
"11101000000000000000100000000000",	-- 1190: 	mulf	%f1, %f0, %f0
"00010100000000100000000000000000",	-- 1191: 	llif	%f2, 1.000000
"00010000000000100011111110000000",	-- 1192: 	lhif	%f2, 1.000000
"00010100000000111010101010011111",	-- 1193: 	llif	%f3, -0.333333
"00010000000000111011111010101010",	-- 1194: 	lhif	%f3, -0.333333
"00010100000001001100110011001101",	-- 1195: 	llif	%f4, 0.200000
"00010000000001000011111001001100",	-- 1196: 	lhif	%f4, 0.200000
"00010100000001010100100100011011",	-- 1197: 	llif	%f5, 0.142857
"00010000000001010011111000010010",	-- 1198: 	lhif	%f5, 0.142857
"11101000001001010010100000000000",	-- 1199: 	mulf	%f5, %f1, %f5
"11100000100001010010000000000000",	-- 1200: 	addf	%f4, %f4, %f5
"11101000001001000010000000000000",	-- 1201: 	mulf	%f4, %f1, %f4
"11100000011001000001100000000000",	-- 1202: 	addf	%f3, %f3, %f4
"11101000001000110000100000000000",	-- 1203: 	mulf	%f1, %f1, %f3
"11100000010000010000100000000000",	-- 1204: 	addf	%f1, %f2, %f1
"11101000000000010000000000000000",	-- 1205: 	mulf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 1206: 	jr	%ra
	-- bgtf_else.8934:
"00010100000000000000000000000000",	-- 1207: 	llif	%f0, -1.000000
"00010000000000001011111110000000",	-- 1208: 	lhif	%f0, -1.000000
"00010100000000010000000000000000",	-- 1209: 	llif	%f1, 1.000000
"00010000000000010011111110000000",	-- 1210: 	lhif	%f1, 1.000000
"10010011110000100000000000000000",	-- 1211: 	lf	%f2, [%sp + 0]
"11101000010000100001100000000000",	-- 1212: 	mulf	%f3, %f2, %f2
"11100000001000110000100000000000",	-- 1213: 	addf	%f1, %f1, %f3
"10110000000111100000000000000001",	-- 1214: 	sf	%f0, [%sp + 1]
"00001100001000000000000000000000",	-- 1215: 	movf	%f0, %f1
"00111111111111100000000000000010",	-- 1216: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1217: 	addi	%sp, %sp, 3
"01011000000000000010101000101110",	-- 1218: 	jal	yj_sqrt
"10101011110111100000000000000011",	-- 1219: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1220: 	lw	%ra, [%sp + 2]
"10010011110000010000000000000001",	-- 1221: 	lf	%f1, [%sp + 1]
"11100000001000000000000000000000",	-- 1222: 	addf	%f0, %f1, %f0
"10010011110000010000000000000000",	-- 1223: 	lf	%f1, [%sp + 0]
"11101100000000010000000000000000",	-- 1224: 	divf	%f0, %f0, %f1
"00010100000000010000000000000000",	-- 1225: 	llif	%f1, 2.000000
"00010000000000010100000000000000",	-- 1226: 	lhif	%f1, 2.000000
"10110000001111100000000000000010",	-- 1227: 	sf	%f1, [%sp + 2]
"00111111111111100000000000000011",	-- 1228: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 1229: 	addi	%sp, %sp, 4
"01011000000000000000010010011100",	-- 1230: 	jal	atan.2520
"10101011110111100000000000000100",	-- 1231: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 1232: 	lw	%ra, [%sp + 3]
"10010011110000010000000000000010",	-- 1233: 	lf	%f1, [%sp + 2]
"11101000001000000000000000000000",	-- 1234: 	mulf	%f0, %f1, %f0
"01001111111000000000000000000000",	-- 1235: 	jr	%ra
	-- fispos.2522:
"00010100000000010000000000000000",	-- 1236: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 1237: 	lhif	%f1, 0.000000
"00100000000000010000000000000011",	-- 1238: 	bgtf	%f0, %f1, bgtf_else.8935
"11001100000000010000000000000000",	-- 1239: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 1240: 	jr	%ra
	-- bgtf_else.8935:
"11001100000000010000000000000001",	-- 1241: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 1242: 	jr	%ra
	-- fisneg.2524:
"00010100000000010000000000000000",	-- 1243: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 1244: 	lhif	%f1, 0.000000
"00100000001000000000000000000011",	-- 1245: 	bgtf	%f1, %f0, bgtf_else.8936
"11001100000000010000000000000000",	-- 1246: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 1247: 	jr	%ra
	-- bgtf_else.8936:
"11001100000000010000000000000001",	-- 1248: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 1249: 	jr	%ra
	-- fiszero.2526:
"00010100000000010000000000000000",	-- 1250: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 1251: 	lhif	%f1, 0.000000
"01011100000000010000000000000000",	-- 1252: 	movf2i	%r1, %f0
"01011100001000100000000000000000",	-- 1253: 	movf2i	%r2, %f1
"00101000001000100000000000000011",	-- 1254: 	bneq	%r1, %r2, bneq_else.8937
"11001100000000010000000000000001",	-- 1255: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 1256: 	jr	%ra
	-- bneq_else.8937:
"11001100000000010000000000000000",	-- 1257: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 1258: 	jr	%ra
	-- fhalf.2528:
"00010100000000010000000000000000",	-- 1259: 	llif	%f1, 0.500000
"00010000000000010011111100000000",	-- 1260: 	lhif	%f1, 0.500000
"11101000000000010000000000000000",	-- 1261: 	mulf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 1262: 	jr	%ra
	-- fsqr.2530:
"11101000000000000000000000000000",	-- 1263: 	mulf	%f0, %f0, %f0
"01001111111000000000000000000000",	-- 1264: 	jr	%ra
	-- fless.2532:
"00100000001000000000000000000011",	-- 1265: 	bgtf	%f1, %f0, bgtf_else.8938
"11001100000000010000000000000000",	-- 1266: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 1267: 	jr	%ra
	-- bgtf_else.8938:
"11001100000000010000000000000001",	-- 1268: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 1269: 	jr	%ra
	-- xor.2565:
"11001100000000110000000000000000",	-- 1270: 	lli	%r3, 0
"00101000001000110000000000000011",	-- 1271: 	bneq	%r1, %r3, bneq_else.8939
"10000100000000100000100000000000",	-- 1272: 	add	%r1, %r0, %r2
"01001111111000000000000000000000",	-- 1273: 	jr	%ra
	-- bneq_else.8939:
"11001100000000010000000000000000",	-- 1274: 	lli	%r1, 0
"00101000010000010000000000000011",	-- 1275: 	bneq	%r2, %r1, bneq_else.8940
"11001100000000010000000000000001",	-- 1276: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 1277: 	jr	%ra
	-- bneq_else.8940:
"11001100000000010000000000000000",	-- 1278: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 1279: 	jr	%ra
	-- sgn.2568:
"10110000000111100000000000000000",	-- 1280: 	sf	%f0, [%sp + 0]
"00111111111111100000000000000001",	-- 1281: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 1282: 	addi	%sp, %sp, 2
"01011000000000000000010011100010",	-- 1283: 	jal	fiszero.2526
"10101011110111100000000000000010",	-- 1284: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 1285: 	lw	%ra, [%sp + 1]
"11001100000000100000000000000000",	-- 1286: 	lli	%r2, 0
"00101000001000100000000000001111",	-- 1287: 	bneq	%r1, %r2, bneq_else.8941
"10010011110000000000000000000000",	-- 1288: 	lf	%f0, [%sp + 0]
"00111111111111100000000000000001",	-- 1289: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 1290: 	addi	%sp, %sp, 2
"01011000000000000000010011010100",	-- 1291: 	jal	fispos.2522
"10101011110111100000000000000010",	-- 1292: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 1293: 	lw	%ra, [%sp + 1]
"11001100000000100000000000000000",	-- 1294: 	lli	%r2, 0
"00101000001000100000000000000100",	-- 1295: 	bneq	%r1, %r2, bneq_else.8942
"00010100000000000000000000000000",	-- 1296: 	llif	%f0, -1.000000
"00010000000000001011111110000000",	-- 1297: 	lhif	%f0, -1.000000
"01001111111000000000000000000000",	-- 1298: 	jr	%ra
	-- bneq_else.8942:
"00010100000000000000000000000000",	-- 1299: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 1300: 	lhif	%f0, 1.000000
"01001111111000000000000000000000",	-- 1301: 	jr	%ra
	-- bneq_else.8941:
"00010100000000000000000000000000",	-- 1302: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 1303: 	lhif	%f0, 0.000000
"01001111111000000000000000000000",	-- 1304: 	jr	%ra
	-- fneg_cond.2570:
"11001100000000100000000000000000",	-- 1305: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 1306: 	bneq	%r1, %r2, bneq_else.8943
"01010100000000000010101001001111",	-- 1307: 	j	yj_fneg
	-- bneq_else.8943:
"01001111111000000000000000000000",	-- 1308: 	jr	%ra
	-- add_mod5.2573:
"10000100001000100000100000000000",	-- 1309: 	add	%r1, %r1, %r2
"11001100000000100000000000000101",	-- 1310: 	lli	%r2, 5
"00110000010000010000000000000100",	-- 1311: 	bgt	%r2, %r1, bgt_else.8944
"11001100000000100000000000000101",	-- 1312: 	lli	%r2, 5
"10001000001000100000100000000000",	-- 1313: 	sub	%r1, %r1, %r2
"01001111111000000000000000000000",	-- 1314: 	jr	%ra
	-- bgt_else.8944:
"01001111111000000000000000000000",	-- 1315: 	jr	%ra
	-- vecset.2576:
"11001100000000100000000000000000",	-- 1316: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 1317: 	add	%r2, %r1, %r2
"10110000000000100000000000000000",	-- 1318: 	sf	%f0, [%r2 + 0]
"11001100000000100000000000000001",	-- 1319: 	lli	%r2, 1
"10000100001000100001000000000000",	-- 1320: 	add	%r2, %r1, %r2
"10110000001000100000000000000000",	-- 1321: 	sf	%f1, [%r2 + 0]
"11001100000000100000000000000010",	-- 1322: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1323: 	add	%r1, %r1, %r2
"10110000010000010000000000000000",	-- 1324: 	sf	%f2, [%r1 + 0]
"01001111111000000000000000000000",	-- 1325: 	jr	%ra
	-- vecfill.2581:
"11001100000000100000000000000000",	-- 1326: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 1327: 	add	%r2, %r1, %r2
"10110000000000100000000000000000",	-- 1328: 	sf	%f0, [%r2 + 0]
"11001100000000100000000000000001",	-- 1329: 	lli	%r2, 1
"10000100001000100001000000000000",	-- 1330: 	add	%r2, %r1, %r2
"10110000000000100000000000000000",	-- 1331: 	sf	%f0, [%r2 + 0]
"11001100000000100000000000000010",	-- 1332: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1333: 	add	%r1, %r1, %r2
"10110000000000010000000000000000",	-- 1334: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1335: 	jr	%ra
	-- vecbzero.2584:
"00010100000000000000000000000000",	-- 1336: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 1337: 	lhif	%f0, 0.000000
"01010100000000000000010100101110",	-- 1338: 	j	vecfill.2581
	-- veccpy.2586:
"11001100000000110000000000000000",	-- 1339: 	lli	%r3, 0
"11001100000001000000000000000000",	-- 1340: 	lli	%r4, 0
"10000100010001000010000000000000",	-- 1341: 	add	%r4, %r2, %r4
"10010000100000000000000000000000",	-- 1342: 	lf	%f0, [%r4 + 0]
"10000100001000110001100000000000",	-- 1343: 	add	%r3, %r1, %r3
"10110000000000110000000000000000",	-- 1344: 	sf	%f0, [%r3 + 0]
"11001100000000110000000000000001",	-- 1345: 	lli	%r3, 1
"11001100000001000000000000000001",	-- 1346: 	lli	%r4, 1
"10000100010001000010000000000000",	-- 1347: 	add	%r4, %r2, %r4
"10010000100000000000000000000000",	-- 1348: 	lf	%f0, [%r4 + 0]
"10000100001000110001100000000000",	-- 1349: 	add	%r3, %r1, %r3
"10110000000000110000000000000000",	-- 1350: 	sf	%f0, [%r3 + 0]
"11001100000000110000000000000010",	-- 1351: 	lli	%r3, 2
"11001100000001000000000000000010",	-- 1352: 	lli	%r4, 2
"10000100010001000001000000000000",	-- 1353: 	add	%r2, %r2, %r4
"10010000010000000000000000000000",	-- 1354: 	lf	%f0, [%r2 + 0]
"10000100001000110000100000000000",	-- 1355: 	add	%r1, %r1, %r3
"10110000000000010000000000000000",	-- 1356: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1357: 	jr	%ra
	-- vecunit_sgn.2594:
"11001100000000110000000000000000",	-- 1358: 	lli	%r3, 0
"10000100001000110001100000000000",	-- 1359: 	add	%r3, %r1, %r3
"10010000011000000000000000000000",	-- 1360: 	lf	%f0, [%r3 + 0]
"00111100010111100000000000000000",	-- 1361: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 1362: 	sw	%r1, [%sp + 1]
"00111111111111100000000000000010",	-- 1363: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1364: 	addi	%sp, %sp, 3
"01011000000000000000010011101111",	-- 1365: 	jal	fsqr.2530
"10101011110111100000000000000011",	-- 1366: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1367: 	lw	%ra, [%sp + 2]
"11001100000000010000000000000001",	-- 1368: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 1369: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 1370: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 1371: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000010",	-- 1372: 	sf	%f0, [%sp + 2]
"00001100001000000000000000000000",	-- 1373: 	movf	%f0, %f1
"00111111111111100000000000000011",	-- 1374: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 1375: 	addi	%sp, %sp, 4
"01011000000000000000010011101111",	-- 1376: 	jal	fsqr.2530
"10101011110111100000000000000100",	-- 1377: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 1378: 	lw	%ra, [%sp + 3]
"10010011110000010000000000000010",	-- 1379: 	lf	%f1, [%sp + 2]
"11100000001000000000000000000000",	-- 1380: 	addf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 1381: 	lli	%r1, 2
"00111011110000100000000000000001",	-- 1382: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 1383: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 1384: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000011",	-- 1385: 	sf	%f0, [%sp + 3]
"00001100001000000000000000000000",	-- 1386: 	movf	%f0, %f1
"00111111111111100000000000000100",	-- 1387: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 1388: 	addi	%sp, %sp, 5
"01011000000000000000010011101111",	-- 1389: 	jal	fsqr.2530
"10101011110111100000000000000101",	-- 1390: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 1391: 	lw	%ra, [%sp + 4]
"10010011110000010000000000000011",	-- 1392: 	lf	%f1, [%sp + 3]
"11100000001000000000000000000000",	-- 1393: 	addf	%f0, %f1, %f0
"00111111111111100000000000000100",	-- 1394: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 1395: 	addi	%sp, %sp, 5
"01011000000000000010101000101110",	-- 1396: 	jal	yj_sqrt
"10101011110111100000000000000101",	-- 1397: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 1398: 	lw	%ra, [%sp + 4]
"10110000000111100000000000000100",	-- 1399: 	sf	%f0, [%sp + 4]
"00111111111111100000000000000101",	-- 1400: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 1401: 	addi	%sp, %sp, 6
"01011000000000000000010011100010",	-- 1402: 	jal	fiszero.2526
"10101011110111100000000000000110",	-- 1403: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 1404: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000000",	-- 1405: 	lli	%r2, 0
"00101000001000100000000000001110",	-- 1406: 	bneq	%r1, %r2, bneq_else.8948
"11001100000000010000000000000000",	-- 1407: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 1408: 	lw	%r2, [%sp + 0]
"00101000010000010000000000000110",	-- 1409: 	bneq	%r2, %r1, bneq_else.8950
"00010100000000000000000000000000",	-- 1410: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 1411: 	lhif	%f0, 1.000000
"10010011110000010000000000000100",	-- 1412: 	lf	%f1, [%sp + 4]
"11101100000000010000000000000000",	-- 1413: 	divf	%f0, %f0, %f1
"01010100000000000000010110001011",	-- 1414: 	j	bneq_cont.8951
	-- bneq_else.8950:
"00010100000000000000000000000000",	-- 1415: 	llif	%f0, -1.000000
"00010000000000001011111110000000",	-- 1416: 	lhif	%f0, -1.000000
"10010011110000010000000000000100",	-- 1417: 	lf	%f1, [%sp + 4]
"11101100000000010000000000000000",	-- 1418: 	divf	%f0, %f0, %f1
	-- bneq_cont.8951:
"01010100000000000000010110001110",	-- 1419: 	j	bneq_cont.8949
	-- bneq_else.8948:
"00010100000000000000000000000000",	-- 1420: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 1421: 	lhif	%f0, 1.000000
	-- bneq_cont.8949:
"11001100000000010000000000000000",	-- 1422: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 1423: 	lli	%r2, 0
"00111011110000110000000000000001",	-- 1424: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 1425: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 1426: 	lf	%f1, [%r2 + 0]
"11101000001000000000100000000000",	-- 1427: 	mulf	%f1, %f1, %f0
"10000100011000010000100000000000",	-- 1428: 	add	%r1, %r3, %r1
"10110000001000010000000000000000",	-- 1429: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000001",	-- 1430: 	lli	%r1, 1
"11001100000000100000000000000001",	-- 1431: 	lli	%r2, 1
"10000100011000100001000000000000",	-- 1432: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 1433: 	lf	%f1, [%r2 + 0]
"11101000001000000000100000000000",	-- 1434: 	mulf	%f1, %f1, %f0
"10000100011000010000100000000000",	-- 1435: 	add	%r1, %r3, %r1
"10110000001000010000000000000000",	-- 1436: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 1437: 	lli	%r1, 2
"11001100000000100000000000000010",	-- 1438: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 1439: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 1440: 	lf	%f1, [%r2 + 0]
"11101000001000000000000000000000",	-- 1441: 	mulf	%f0, %f1, %f0
"10000100011000010000100000000000",	-- 1442: 	add	%r1, %r3, %r1
"10110000000000010000000000000000",	-- 1443: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1444: 	jr	%ra
	-- veciprod.2597:
"11001100000000110000000000000000",	-- 1445: 	lli	%r3, 0
"10000100001000110001100000000000",	-- 1446: 	add	%r3, %r1, %r3
"10010000011000000000000000000000",	-- 1447: 	lf	%f0, [%r3 + 0]
"11001100000000110000000000000000",	-- 1448: 	lli	%r3, 0
"10000100010000110001100000000000",	-- 1449: 	add	%r3, %r2, %r3
"10010000011000010000000000000000",	-- 1450: 	lf	%f1, [%r3 + 0]
"11101000000000010000000000000000",	-- 1451: 	mulf	%f0, %f0, %f1
"11001100000000110000000000000001",	-- 1452: 	lli	%r3, 1
"10000100001000110001100000000000",	-- 1453: 	add	%r3, %r1, %r3
"10010000011000010000000000000000",	-- 1454: 	lf	%f1, [%r3 + 0]
"11001100000000110000000000000001",	-- 1455: 	lli	%r3, 1
"10000100010000110001100000000000",	-- 1456: 	add	%r3, %r2, %r3
"10010000011000100000000000000000",	-- 1457: 	lf	%f2, [%r3 + 0]
"11101000001000100000100000000000",	-- 1458: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 1459: 	addf	%f0, %f0, %f1
"11001100000000110000000000000010",	-- 1460: 	lli	%r3, 2
"10000100001000110000100000000000",	-- 1461: 	add	%r1, %r1, %r3
"10010000001000010000000000000000",	-- 1462: 	lf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 1463: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 1464: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 1465: 	lf	%f2, [%r1 + 0]
"11101000001000100000100000000000",	-- 1466: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 1467: 	addf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 1468: 	jr	%ra
	-- veciprod2.2600:
"11001100000000100000000000000000",	-- 1469: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 1470: 	add	%r2, %r1, %r2
"10010000010000110000000000000000",	-- 1471: 	lf	%f3, [%r2 + 0]
"11101000011000000000000000000000",	-- 1472: 	mulf	%f0, %f3, %f0
"11001100000000100000000000000001",	-- 1473: 	lli	%r2, 1
"10000100001000100001000000000000",	-- 1474: 	add	%r2, %r1, %r2
"10010000010000110000000000000000",	-- 1475: 	lf	%f3, [%r2 + 0]
"11101000011000010000100000000000",	-- 1476: 	mulf	%f1, %f3, %f1
"11100000000000010000000000000000",	-- 1477: 	addf	%f0, %f0, %f1
"11001100000000100000000000000010",	-- 1478: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1479: 	add	%r1, %r1, %r2
"10010000001000010000000000000000",	-- 1480: 	lf	%f1, [%r1 + 0]
"11101000001000100000100000000000",	-- 1481: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 1482: 	addf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 1483: 	jr	%ra
	-- vecaccum.2605:
"11001100000000110000000000000000",	-- 1484: 	lli	%r3, 0
"11001100000001000000000000000000",	-- 1485: 	lli	%r4, 0
"10000100001001000010000000000000",	-- 1486: 	add	%r4, %r1, %r4
"10010000100000010000000000000000",	-- 1487: 	lf	%f1, [%r4 + 0]
"11001100000001000000000000000000",	-- 1488: 	lli	%r4, 0
"10000100010001000010000000000000",	-- 1489: 	add	%r4, %r2, %r4
"10010000100000100000000000000000",	-- 1490: 	lf	%f2, [%r4 + 0]
"11101000000000100001000000000000",	-- 1491: 	mulf	%f2, %f0, %f2
"11100000001000100000100000000000",	-- 1492: 	addf	%f1, %f1, %f2
"10000100001000110001100000000000",	-- 1493: 	add	%r3, %r1, %r3
"10110000001000110000000000000000",	-- 1494: 	sf	%f1, [%r3 + 0]
"11001100000000110000000000000001",	-- 1495: 	lli	%r3, 1
"11001100000001000000000000000001",	-- 1496: 	lli	%r4, 1
"10000100001001000010000000000000",	-- 1497: 	add	%r4, %r1, %r4
"10010000100000010000000000000000",	-- 1498: 	lf	%f1, [%r4 + 0]
"11001100000001000000000000000001",	-- 1499: 	lli	%r4, 1
"10000100010001000010000000000000",	-- 1500: 	add	%r4, %r2, %r4
"10010000100000100000000000000000",	-- 1501: 	lf	%f2, [%r4 + 0]
"11101000000000100001000000000000",	-- 1502: 	mulf	%f2, %f0, %f2
"11100000001000100000100000000000",	-- 1503: 	addf	%f1, %f1, %f2
"10000100001000110001100000000000",	-- 1504: 	add	%r3, %r1, %r3
"10110000001000110000000000000000",	-- 1505: 	sf	%f1, [%r3 + 0]
"11001100000000110000000000000010",	-- 1506: 	lli	%r3, 2
"11001100000001000000000000000010",	-- 1507: 	lli	%r4, 2
"10000100001001000010000000000000",	-- 1508: 	add	%r4, %r1, %r4
"10010000100000010000000000000000",	-- 1509: 	lf	%f1, [%r4 + 0]
"11001100000001000000000000000010",	-- 1510: 	lli	%r4, 2
"10000100010001000001000000000000",	-- 1511: 	add	%r2, %r2, %r4
"10010000010000100000000000000000",	-- 1512: 	lf	%f2, [%r2 + 0]
"11101000000000100000000000000000",	-- 1513: 	mulf	%f0, %f0, %f2
"11100000001000000000000000000000",	-- 1514: 	addf	%f0, %f1, %f0
"10000100001000110000100000000000",	-- 1515: 	add	%r1, %r1, %r3
"10110000000000010000000000000000",	-- 1516: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1517: 	jr	%ra
	-- vecadd.2609:
"11001100000000110000000000000000",	-- 1518: 	lli	%r3, 0
"11001100000001000000000000000000",	-- 1519: 	lli	%r4, 0
"10000100001001000010000000000000",	-- 1520: 	add	%r4, %r1, %r4
"10010000100000000000000000000000",	-- 1521: 	lf	%f0, [%r4 + 0]
"11001100000001000000000000000000",	-- 1522: 	lli	%r4, 0
"10000100010001000010000000000000",	-- 1523: 	add	%r4, %r2, %r4
"10010000100000010000000000000000",	-- 1524: 	lf	%f1, [%r4 + 0]
"11100000000000010000000000000000",	-- 1525: 	addf	%f0, %f0, %f1
"10000100001000110001100000000000",	-- 1526: 	add	%r3, %r1, %r3
"10110000000000110000000000000000",	-- 1527: 	sf	%f0, [%r3 + 0]
"11001100000000110000000000000001",	-- 1528: 	lli	%r3, 1
"11001100000001000000000000000001",	-- 1529: 	lli	%r4, 1
"10000100001001000010000000000000",	-- 1530: 	add	%r4, %r1, %r4
"10010000100000000000000000000000",	-- 1531: 	lf	%f0, [%r4 + 0]
"11001100000001000000000000000001",	-- 1532: 	lli	%r4, 1
"10000100010001000010000000000000",	-- 1533: 	add	%r4, %r2, %r4
"10010000100000010000000000000000",	-- 1534: 	lf	%f1, [%r4 + 0]
"11100000000000010000000000000000",	-- 1535: 	addf	%f0, %f0, %f1
"10000100001000110001100000000000",	-- 1536: 	add	%r3, %r1, %r3
"10110000000000110000000000000000",	-- 1537: 	sf	%f0, [%r3 + 0]
"11001100000000110000000000000010",	-- 1538: 	lli	%r3, 2
"11001100000001000000000000000010",	-- 1539: 	lli	%r4, 2
"10000100001001000010000000000000",	-- 1540: 	add	%r4, %r1, %r4
"10010000100000000000000000000000",	-- 1541: 	lf	%f0, [%r4 + 0]
"11001100000001000000000000000010",	-- 1542: 	lli	%r4, 2
"10000100010001000001000000000000",	-- 1543: 	add	%r2, %r2, %r4
"10010000010000010000000000000000",	-- 1544: 	lf	%f1, [%r2 + 0]
"11100000000000010000000000000000",	-- 1545: 	addf	%f0, %f0, %f1
"10000100001000110000100000000000",	-- 1546: 	add	%r1, %r1, %r3
"10110000000000010000000000000000",	-- 1547: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1548: 	jr	%ra
	-- vecscale.2615:
"11001100000000100000000000000000",	-- 1549: 	lli	%r2, 0
"11001100000000110000000000000000",	-- 1550: 	lli	%r3, 0
"10000100001000110001100000000000",	-- 1551: 	add	%r3, %r1, %r3
"10010000011000010000000000000000",	-- 1552: 	lf	%f1, [%r3 + 0]
"11101000001000000000100000000000",	-- 1553: 	mulf	%f1, %f1, %f0
"10000100001000100001000000000000",	-- 1554: 	add	%r2, %r1, %r2
"10110000001000100000000000000000",	-- 1555: 	sf	%f1, [%r2 + 0]
"11001100000000100000000000000001",	-- 1556: 	lli	%r2, 1
"11001100000000110000000000000001",	-- 1557: 	lli	%r3, 1
"10000100001000110001100000000000",	-- 1558: 	add	%r3, %r1, %r3
"10010000011000010000000000000000",	-- 1559: 	lf	%f1, [%r3 + 0]
"11101000001000000000100000000000",	-- 1560: 	mulf	%f1, %f1, %f0
"10000100001000100001000000000000",	-- 1561: 	add	%r2, %r1, %r2
"10110000001000100000000000000000",	-- 1562: 	sf	%f1, [%r2 + 0]
"11001100000000100000000000000010",	-- 1563: 	lli	%r2, 2
"11001100000000110000000000000010",	-- 1564: 	lli	%r3, 2
"10000100001000110001100000000000",	-- 1565: 	add	%r3, %r1, %r3
"10010000011000010000000000000000",	-- 1566: 	lf	%f1, [%r3 + 0]
"11101000001000000000000000000000",	-- 1567: 	mulf	%f0, %f1, %f0
"10000100001000100000100000000000",	-- 1568: 	add	%r1, %r1, %r2
"10110000000000010000000000000000",	-- 1569: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1570: 	jr	%ra
	-- vecaccumv.2618:
"11001100000001000000000000000000",	-- 1571: 	lli	%r4, 0
"11001100000001010000000000000000",	-- 1572: 	lli	%r5, 0
"10000100001001010010100000000000",	-- 1573: 	add	%r5, %r1, %r5
"10010000101000000000000000000000",	-- 1574: 	lf	%f0, [%r5 + 0]
"11001100000001010000000000000000",	-- 1575: 	lli	%r5, 0
"10000100010001010010100000000000",	-- 1576: 	add	%r5, %r2, %r5
"10010000101000010000000000000000",	-- 1577: 	lf	%f1, [%r5 + 0]
"11001100000001010000000000000000",	-- 1578: 	lli	%r5, 0
"10000100011001010010100000000000",	-- 1579: 	add	%r5, %r3, %r5
"10010000101000100000000000000000",	-- 1580: 	lf	%f2, [%r5 + 0]
"11101000001000100000100000000000",	-- 1581: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 1582: 	addf	%f0, %f0, %f1
"10000100001001000010000000000000",	-- 1583: 	add	%r4, %r1, %r4
"10110000000001000000000000000000",	-- 1584: 	sf	%f0, [%r4 + 0]
"11001100000001000000000000000001",	-- 1585: 	lli	%r4, 1
"11001100000001010000000000000001",	-- 1586: 	lli	%r5, 1
"10000100001001010010100000000000",	-- 1587: 	add	%r5, %r1, %r5
"10010000101000000000000000000000",	-- 1588: 	lf	%f0, [%r5 + 0]
"11001100000001010000000000000001",	-- 1589: 	lli	%r5, 1
"10000100010001010010100000000000",	-- 1590: 	add	%r5, %r2, %r5
"10010000101000010000000000000000",	-- 1591: 	lf	%f1, [%r5 + 0]
"11001100000001010000000000000001",	-- 1592: 	lli	%r5, 1
"10000100011001010010100000000000",	-- 1593: 	add	%r5, %r3, %r5
"10010000101000100000000000000000",	-- 1594: 	lf	%f2, [%r5 + 0]
"11101000001000100000100000000000",	-- 1595: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 1596: 	addf	%f0, %f0, %f1
"10000100001001000010000000000000",	-- 1597: 	add	%r4, %r1, %r4
"10110000000001000000000000000000",	-- 1598: 	sf	%f0, [%r4 + 0]
"11001100000001000000000000000010",	-- 1599: 	lli	%r4, 2
"11001100000001010000000000000010",	-- 1600: 	lli	%r5, 2
"10000100001001010010100000000000",	-- 1601: 	add	%r5, %r1, %r5
"10010000101000000000000000000000",	-- 1602: 	lf	%f0, [%r5 + 0]
"11001100000001010000000000000010",	-- 1603: 	lli	%r5, 2
"10000100010001010001000000000000",	-- 1604: 	add	%r2, %r2, %r5
"10010000010000010000000000000000",	-- 1605: 	lf	%f1, [%r2 + 0]
"11001100000000100000000000000010",	-- 1606: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 1607: 	add	%r2, %r3, %r2
"10010000010000100000000000000000",	-- 1608: 	lf	%f2, [%r2 + 0]
"11101000001000100000100000000000",	-- 1609: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 1610: 	addf	%f0, %f0, %f1
"10000100001001000000100000000000",	-- 1611: 	add	%r1, %r1, %r4
"10110000000000010000000000000000",	-- 1612: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1613: 	jr	%ra
	-- o_texturetype.2622:
"00111000001000010000000000000000",	-- 1614: 	lw	%r1, [%r1 + 0]
"01001111111000000000000000000000",	-- 1615: 	jr	%ra
	-- o_form.2624:
"00111000001000010000000000000001",	-- 1616: 	lw	%r1, [%r1 + 1]
"01001111111000000000000000000000",	-- 1617: 	jr	%ra
	-- o_reflectiontype.2626:
"00111000001000010000000000000010",	-- 1618: 	lw	%r1, [%r1 + 2]
"01001111111000000000000000000000",	-- 1619: 	jr	%ra
	-- o_isinvert.2628:
"00111000001000010000000000000110",	-- 1620: 	lw	%r1, [%r1 + 6]
"01001111111000000000000000000000",	-- 1621: 	jr	%ra
	-- o_isrot.2630:
"00111000001000010000000000000011",	-- 1622: 	lw	%r1, [%r1 + 3]
"01001111111000000000000000000000",	-- 1623: 	jr	%ra
	-- o_param_a.2632:
"00111000001000010000000000000100",	-- 1624: 	lw	%r1, [%r1 + 4]
"11001100000000100000000000000000",	-- 1625: 	lli	%r2, 0
"10000100001000100000100000000000",	-- 1626: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1627: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1628: 	jr	%ra
	-- o_param_b.2634:
"00111000001000010000000000000100",	-- 1629: 	lw	%r1, [%r1 + 4]
"11001100000000100000000000000001",	-- 1630: 	lli	%r2, 1
"10000100001000100000100000000000",	-- 1631: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1632: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1633: 	jr	%ra
	-- o_param_c.2636:
"00111000001000010000000000000100",	-- 1634: 	lw	%r1, [%r1 + 4]
"11001100000000100000000000000010",	-- 1635: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1636: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1637: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1638: 	jr	%ra
	-- o_param_abc.2638:
"00111000001000010000000000000100",	-- 1639: 	lw	%r1, [%r1 + 4]
"01001111111000000000000000000000",	-- 1640: 	jr	%ra
	-- o_param_x.2640:
"00111000001000010000000000000101",	-- 1641: 	lw	%r1, [%r1 + 5]
"11001100000000100000000000000000",	-- 1642: 	lli	%r2, 0
"10000100001000100000100000000000",	-- 1643: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1644: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1645: 	jr	%ra
	-- o_param_y.2642:
"00111000001000010000000000000101",	-- 1646: 	lw	%r1, [%r1 + 5]
"11001100000000100000000000000001",	-- 1647: 	lli	%r2, 1
"10000100001000100000100000000000",	-- 1648: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1649: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1650: 	jr	%ra
	-- o_param_z.2644:
"00111000001000010000000000000101",	-- 1651: 	lw	%r1, [%r1 + 5]
"11001100000000100000000000000010",	-- 1652: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1653: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1654: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1655: 	jr	%ra
	-- o_diffuse.2646:
"00111000001000010000000000000111",	-- 1656: 	lw	%r1, [%r1 + 7]
"11001100000000100000000000000000",	-- 1657: 	lli	%r2, 0
"10000100001000100000100000000000",	-- 1658: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1659: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1660: 	jr	%ra
	-- o_hilight.2648:
"00111000001000010000000000000111",	-- 1661: 	lw	%r1, [%r1 + 7]
"11001100000000100000000000000001",	-- 1662: 	lli	%r2, 1
"10000100001000100000100000000000",	-- 1663: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1664: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1665: 	jr	%ra
	-- o_color_red.2650:
"00111000001000010000000000001000",	-- 1666: 	lw	%r1, [%r1 + 8]
"11001100000000100000000000000000",	-- 1667: 	lli	%r2, 0
"10000100001000100000100000000000",	-- 1668: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1669: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1670: 	jr	%ra
	-- o_color_green.2652:
"00111000001000010000000000001000",	-- 1671: 	lw	%r1, [%r1 + 8]
"11001100000000100000000000000001",	-- 1672: 	lli	%r2, 1
"10000100001000100000100000000000",	-- 1673: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1674: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1675: 	jr	%ra
	-- o_color_blue.2654:
"00111000001000010000000000001000",	-- 1676: 	lw	%r1, [%r1 + 8]
"11001100000000100000000000000010",	-- 1677: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1678: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1679: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1680: 	jr	%ra
	-- o_param_r1.2656:
"00111000001000010000000000001001",	-- 1681: 	lw	%r1, [%r1 + 9]
"11001100000000100000000000000000",	-- 1682: 	lli	%r2, 0
"10000100001000100000100000000000",	-- 1683: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1684: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1685: 	jr	%ra
	-- o_param_r2.2658:
"00111000001000010000000000001001",	-- 1686: 	lw	%r1, [%r1 + 9]
"11001100000000100000000000000001",	-- 1687: 	lli	%r2, 1
"10000100001000100000100000000000",	-- 1688: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1689: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1690: 	jr	%ra
	-- o_param_r3.2660:
"00111000001000010000000000001001",	-- 1691: 	lw	%r1, [%r1 + 9]
"11001100000000100000000000000010",	-- 1692: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1693: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1694: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1695: 	jr	%ra
	-- o_param_ctbl.2662:
"00111000001000010000000000001010",	-- 1696: 	lw	%r1, [%r1 + 10]
"01001111111000000000000000000000",	-- 1697: 	jr	%ra
	-- p_rgb.2664:
"00111000001000010000000000000000",	-- 1698: 	lw	%r1, [%r1 + 0]
"01001111111000000000000000000000",	-- 1699: 	jr	%ra
	-- p_intersection_points.2666:
"00111000001000010000000000000001",	-- 1700: 	lw	%r1, [%r1 + 1]
"01001111111000000000000000000000",	-- 1701: 	jr	%ra
	-- p_surface_ids.2668:
"00111000001000010000000000000010",	-- 1702: 	lw	%r1, [%r1 + 2]
"01001111111000000000000000000000",	-- 1703: 	jr	%ra
	-- p_calc_diffuse.2670:
"00111000001000010000000000000011",	-- 1704: 	lw	%r1, [%r1 + 3]
"01001111111000000000000000000000",	-- 1705: 	jr	%ra
	-- p_energy.2672:
"00111000001000010000000000000100",	-- 1706: 	lw	%r1, [%r1 + 4]
"01001111111000000000000000000000",	-- 1707: 	jr	%ra
	-- p_received_ray_20percent.2674:
"00111000001000010000000000000101",	-- 1708: 	lw	%r1, [%r1 + 5]
"01001111111000000000000000000000",	-- 1709: 	jr	%ra
	-- p_group_id.2676:
"00111000001000010000000000000110",	-- 1710: 	lw	%r1, [%r1 + 6]
"11001100000000100000000000000000",	-- 1711: 	lli	%r2, 0
"10000100001000100000100000000000",	-- 1712: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 1713: 	lw	%r1, [%r1 + 0]
"01001111111000000000000000000000",	-- 1714: 	jr	%ra
	-- p_set_group_id.2678:
"00111000001000010000000000000110",	-- 1715: 	lw	%r1, [%r1 + 6]
"11001100000000110000000000000000",	-- 1716: 	lli	%r3, 0
"10000100001000110000100000000000",	-- 1717: 	add	%r1, %r1, %r3
"00111100010000010000000000000000",	-- 1718: 	sw	%r2, [%r1 + 0]
"01001111111000000000000000000000",	-- 1719: 	jr	%ra
	-- p_nvectors.2681:
"00111000001000010000000000000111",	-- 1720: 	lw	%r1, [%r1 + 7]
"01001111111000000000000000000000",	-- 1721: 	jr	%ra
	-- d_vec.2683:
"00111000001000010000000000000000",	-- 1722: 	lw	%r1, [%r1 + 0]
"01001111111000000000000000000000",	-- 1723: 	jr	%ra
	-- d_const.2685:
"00111000001000010000000000000001",	-- 1724: 	lw	%r1, [%r1 + 1]
"01001111111000000000000000000000",	-- 1725: 	jr	%ra
	-- r_surface_id.2687:
"00111000001000010000000000000000",	-- 1726: 	lw	%r1, [%r1 + 0]
"01001111111000000000000000000000",	-- 1727: 	jr	%ra
	-- r_dvec.2689:
"00111000001000010000000000000001",	-- 1728: 	lw	%r1, [%r1 + 1]
"01001111111000000000000000000000",	-- 1729: 	jr	%ra
	-- r_bright.2691:
"10010000001000000000000000000010",	-- 1730: 	lf	%f0, [%r1 + 2]
"01001111111000000000000000000000",	-- 1731: 	jr	%ra
	-- rad.2693:
"00010100000000011111100110011000",	-- 1732: 	llif	%f1, 0.017453
"00010000000000010011110010001110",	-- 1733: 	lhif	%f1, 0.017453
"11101000000000010000000000000000",	-- 1734: 	mulf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 1735: 	jr	%ra
	-- read_screen_settings.2695:
"00111011011000010000000000000101",	-- 1736: 	lw	%r1, [%r27 + 5]
"00111011011000100000000000000100",	-- 1737: 	lw	%r2, [%r27 + 4]
"00111011011000110000000000000011",	-- 1738: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 1739: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 1740: 	lw	%r5, [%r27 + 1]
"11001100000001100000000000000000",	-- 1741: 	lli	%r6, 0
"00111100001111100000000000000000",	-- 1742: 	sw	%r1, [%sp + 0]
"00111100011111100000000000000001",	-- 1743: 	sw	%r3, [%sp + 1]
"00111100100111100000000000000010",	-- 1744: 	sw	%r4, [%sp + 2]
"00111100010111100000000000000011",	-- 1745: 	sw	%r2, [%sp + 3]
"00111100110111100000000000000100",	-- 1746: 	sw	%r6, [%sp + 4]
"00111100101111100000000000000101",	-- 1747: 	sw	%r5, [%sp + 5]
"00111111111111100000000000000110",	-- 1748: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 1749: 	addi	%sp, %sp, 7
"01011000000000000010101000111111",	-- 1750: 	jal	yj_read_float
"10101011110111100000000000000111",	-- 1751: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 1752: 	lw	%ra, [%sp + 6]
"00111011110000010000000000000100",	-- 1753: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000101",	-- 1754: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 1755: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1756: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 1757: 	lli	%r1, 1
"00111100001111100000000000000110",	-- 1758: 	sw	%r1, [%sp + 6]
"00111111111111100000000000000111",	-- 1759: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 1760: 	addi	%sp, %sp, 8
"01011000000000000010101000111111",	-- 1761: 	jal	yj_read_float
"10101011110111100000000000001000",	-- 1762: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 1763: 	lw	%ra, [%sp + 7]
"00111011110000010000000000000110",	-- 1764: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000101",	-- 1765: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 1766: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1767: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 1768: 	lli	%r1, 2
"00111100001111100000000000000111",	-- 1769: 	sw	%r1, [%sp + 7]
"00111111111111100000000000001000",	-- 1770: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 1771: 	addi	%sp, %sp, 9
"01011000000000000010101000111111",	-- 1772: 	jal	yj_read_float
"10101011110111100000000000001001",	-- 1773: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 1774: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000111",	-- 1775: 	lw	%r1, [%sp + 7]
"00111011110000100000000000000101",	-- 1776: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 1777: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1778: 	sf	%f0, [%r1 + 0]
"00111111111111100000000000001000",	-- 1779: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 1780: 	addi	%sp, %sp, 9
"01011000000000000010101000111111",	-- 1781: 	jal	yj_read_float
"10101011110111100000000000001001",	-- 1782: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 1783: 	lw	%ra, [%sp + 8]
"00111111111111100000000000001000",	-- 1784: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 1785: 	addi	%sp, %sp, 9
"01011000000000000000011011000100",	-- 1786: 	jal	rad.2693
"10101011110111100000000000001001",	-- 1787: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 1788: 	lw	%ra, [%sp + 8]
"10110000000111100000000000001000",	-- 1789: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 1790: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 1791: 	addi	%sp, %sp, 10
"01011000000000000000010010010110",	-- 1792: 	jal	cos.2518
"10101011110111100000000000001010",	-- 1793: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 1794: 	lw	%ra, [%sp + 9]
"10010011110000010000000000001000",	-- 1795: 	lf	%f1, [%sp + 8]
"10110000000111100000000000001001",	-- 1796: 	sf	%f0, [%sp + 9]
"00001100001000000000000000000000",	-- 1797: 	movf	%f0, %f1
"00111111111111100000000000001010",	-- 1798: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 1799: 	addi	%sp, %sp, 11
"01011000000000000000010001010111",	-- 1800: 	jal	sin.2516
"10101011110111100000000000001011",	-- 1801: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 1802: 	lw	%ra, [%sp + 10]
"10110000000111100000000000001010",	-- 1803: 	sf	%f0, [%sp + 10]
"00111111111111100000000000001011",	-- 1804: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 1805: 	addi	%sp, %sp, 12
"01011000000000000010101000111111",	-- 1806: 	jal	yj_read_float
"10101011110111100000000000001100",	-- 1807: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 1808: 	lw	%ra, [%sp + 11]
"00111111111111100000000000001011",	-- 1809: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 1810: 	addi	%sp, %sp, 12
"01011000000000000000011011000100",	-- 1811: 	jal	rad.2693
"10101011110111100000000000001100",	-- 1812: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 1813: 	lw	%ra, [%sp + 11]
"10110000000111100000000000001011",	-- 1814: 	sf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 1815: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 1816: 	addi	%sp, %sp, 13
"01011000000000000000010010010110",	-- 1817: 	jal	cos.2518
"10101011110111100000000000001101",	-- 1818: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 1819: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001011",	-- 1820: 	lf	%f1, [%sp + 11]
"10110000000111100000000000001100",	-- 1821: 	sf	%f0, [%sp + 12]
"00001100001000000000000000000000",	-- 1822: 	movf	%f0, %f1
"00111111111111100000000000001101",	-- 1823: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 1824: 	addi	%sp, %sp, 14
"01011000000000000000010001010111",	-- 1825: 	jal	sin.2516
"10101011110111100000000000001110",	-- 1826: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 1827: 	lw	%ra, [%sp + 13]
"11001100000000010000000000000000",	-- 1828: 	lli	%r1, 0
"10010011110000010000000000001001",	-- 1829: 	lf	%f1, [%sp + 9]
"11101000001000000001000000000000",	-- 1830: 	mulf	%f2, %f1, %f0
"00010100000000110000000000000000",	-- 1831: 	llif	%f3, 200.000000
"00010000000000110100001101001000",	-- 1832: 	lhif	%f3, 200.000000
"11101000010000110001000000000000",	-- 1833: 	mulf	%f2, %f2, %f3
"00111011110000100000000000000011",	-- 1834: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 1835: 	add	%r1, %r2, %r1
"10110000010000010000000000000000",	-- 1836: 	sf	%f2, [%r1 + 0]
"11001100000000010000000000000001",	-- 1837: 	lli	%r1, 1
"00010100000000100000000000000000",	-- 1838: 	llif	%f2, -200.000000
"00010000000000101100001101001000",	-- 1839: 	lhif	%f2, -200.000000
"10010011110000110000000000001010",	-- 1840: 	lf	%f3, [%sp + 10]
"11101000011000100001000000000000",	-- 1841: 	mulf	%f2, %f3, %f2
"10000100010000010000100000000000",	-- 1842: 	add	%r1, %r2, %r1
"10110000010000010000000000000000",	-- 1843: 	sf	%f2, [%r1 + 0]
"11001100000000010000000000000010",	-- 1844: 	lli	%r1, 2
"10010011110000100000000000001100",	-- 1845: 	lf	%f2, [%sp + 12]
"11101000001000100010000000000000",	-- 1846: 	mulf	%f4, %f1, %f2
"00010100000001010000000000000000",	-- 1847: 	llif	%f5, 200.000000
"00010000000001010100001101001000",	-- 1848: 	lhif	%f5, 200.000000
"11101000100001010010000000000000",	-- 1849: 	mulf	%f4, %f4, %f5
"10000100010000010000100000000000",	-- 1850: 	add	%r1, %r2, %r1
"10110000100000010000000000000000",	-- 1851: 	sf	%f4, [%r1 + 0]
"11001100000000010000000000000000",	-- 1852: 	lli	%r1, 0
"00111011110000110000000000000010",	-- 1853: 	lw	%r3, [%sp + 2]
"10000100011000010000100000000000",	-- 1854: 	add	%r1, %r3, %r1
"10110000010000010000000000000000",	-- 1855: 	sf	%f2, [%r1 + 0]
"11001100000000010000000000000001",	-- 1856: 	lli	%r1, 1
"00010100000001000000000000000000",	-- 1857: 	llif	%f4, 0.000000
"00010000000001000000000000000000",	-- 1858: 	lhif	%f4, 0.000000
"10000100011000010000100000000000",	-- 1859: 	add	%r1, %r3, %r1
"10110000100000010000000000000000",	-- 1860: 	sf	%f4, [%r1 + 0]
"11001100000000010000000000000010",	-- 1861: 	lli	%r1, 2
"10110000000111100000000000001101",	-- 1862: 	sf	%f0, [%sp + 13]
"00111100001111100000000000001110",	-- 1863: 	sw	%r1, [%sp + 14]
"00111111111111100000000000001111",	-- 1864: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 1865: 	addi	%sp, %sp, 16
"01011000000000000010101001001111",	-- 1866: 	jal	yj_fneg
"10101011110111100000000000010000",	-- 1867: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 1868: 	lw	%ra, [%sp + 15]
"00111011110000010000000000001110",	-- 1869: 	lw	%r1, [%sp + 14]
"00111011110000100000000000000010",	-- 1870: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 1871: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1872: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 1873: 	lli	%r1, 0
"10010011110000000000000000001010",	-- 1874: 	lf	%f0, [%sp + 10]
"00111100001111100000000000001111",	-- 1875: 	sw	%r1, [%sp + 15]
"00111111111111100000000000010000",	-- 1876: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 1877: 	addi	%sp, %sp, 17
"01011000000000000010101001001111",	-- 1878: 	jal	yj_fneg
"10101011110111100000000000010001",	-- 1879: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 1880: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001101",	-- 1881: 	lf	%f1, [%sp + 13]
"11101000000000010000000000000000",	-- 1882: 	mulf	%f0, %f0, %f1
"00111011110000010000000000001111",	-- 1883: 	lw	%r1, [%sp + 15]
"00111011110000100000000000000001",	-- 1884: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 1885: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1886: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 1887: 	lli	%r1, 1
"10010011110000000000000000001001",	-- 1888: 	lf	%f0, [%sp + 9]
"00111100001111100000000000010000",	-- 1889: 	sw	%r1, [%sp + 16]
"00111111111111100000000000010001",	-- 1890: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 1891: 	addi	%sp, %sp, 18
"01011000000000000010101001001111",	-- 1892: 	jal	yj_fneg
"10101011110111100000000000010010",	-- 1893: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 1894: 	lw	%ra, [%sp + 17]
"00111011110000010000000000010000",	-- 1895: 	lw	%r1, [%sp + 16]
"00111011110000100000000000000001",	-- 1896: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 1897: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1898: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 1899: 	lli	%r1, 2
"10010011110000000000000000001010",	-- 1900: 	lf	%f0, [%sp + 10]
"00111100001111100000000000010001",	-- 1901: 	sw	%r1, [%sp + 17]
"00111111111111100000000000010010",	-- 1902: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 1903: 	addi	%sp, %sp, 19
"01011000000000000010101001001111",	-- 1904: 	jal	yj_fneg
"10101011110111100000000000010011",	-- 1905: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 1906: 	lw	%ra, [%sp + 18]
"10010011110000010000000000001100",	-- 1907: 	lf	%f1, [%sp + 12]
"11101000000000010000000000000000",	-- 1908: 	mulf	%f0, %f0, %f1
"00111011110000010000000000010001",	-- 1909: 	lw	%r1, [%sp + 17]
"00111011110000100000000000000001",	-- 1910: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 1911: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1912: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 1913: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 1914: 	lli	%r2, 0
"00111011110000110000000000000101",	-- 1915: 	lw	%r3, [%sp + 5]
"10000100011000100001000000000000",	-- 1916: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 1917: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000000",	-- 1918: 	lli	%r2, 0
"00111011110001000000000000000011",	-- 1919: 	lw	%r4, [%sp + 3]
"10000100100000100001000000000000",	-- 1920: 	add	%r2, %r4, %r2
"10010000010000010000000000000000",	-- 1921: 	lf	%f1, [%r2 + 0]
"11100100000000010000000000000000",	-- 1922: 	subf	%f0, %f0, %f1
"00111011110000100000000000000000",	-- 1923: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 1924: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1925: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 1926: 	lli	%r1, 1
"11001100000001010000000000000001",	-- 1927: 	lli	%r5, 1
"10000100011001010010100000000000",	-- 1928: 	add	%r5, %r3, %r5
"10010000101000000000000000000000",	-- 1929: 	lf	%f0, [%r5 + 0]
"11001100000001010000000000000001",	-- 1930: 	lli	%r5, 1
"10000100100001010010100000000000",	-- 1931: 	add	%r5, %r4, %r5
"10010000101000010000000000000000",	-- 1932: 	lf	%f1, [%r5 + 0]
"11100100000000010000000000000000",	-- 1933: 	subf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 1934: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1935: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 1936: 	lli	%r1, 2
"11001100000001010000000000000010",	-- 1937: 	lli	%r5, 2
"10000100011001010001100000000000",	-- 1938: 	add	%r3, %r3, %r5
"10010000011000000000000000000000",	-- 1939: 	lf	%f0, [%r3 + 0]
"11001100000000110000000000000010",	-- 1940: 	lli	%r3, 2
"10000100100000110001100000000000",	-- 1941: 	add	%r3, %r4, %r3
"10010000011000010000000000000000",	-- 1942: 	lf	%f1, [%r3 + 0]
"11100100000000010000000000000000",	-- 1943: 	subf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 1944: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1945: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1946: 	jr	%ra
	-- read_light.2697:
"00111011011000010000000000000010",	-- 1947: 	lw	%r1, [%r27 + 2]
"00111011011000100000000000000001",	-- 1948: 	lw	%r2, [%r27 + 1]
"00111100010111100000000000000000",	-- 1949: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 1950: 	sw	%r1, [%sp + 1]
"00111111111111100000000000000010",	-- 1951: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1952: 	addi	%sp, %sp, 3
"01011000000000000010101000110010",	-- 1953: 	jal	yj_read_int
"10101011110111100000000000000011",	-- 1954: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1955: 	lw	%ra, [%sp + 2]
"00111111111111100000000000000010",	-- 1956: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1957: 	addi	%sp, %sp, 3
"01011000000000000010101000111111",	-- 1958: 	jal	yj_read_float
"10101011110111100000000000000011",	-- 1959: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1960: 	lw	%ra, [%sp + 2]
"00111111111111100000000000000010",	-- 1961: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1962: 	addi	%sp, %sp, 3
"01011000000000000000011011000100",	-- 1963: 	jal	rad.2693
"10101011110111100000000000000011",	-- 1964: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1965: 	lw	%ra, [%sp + 2]
"10110000000111100000000000000010",	-- 1966: 	sf	%f0, [%sp + 2]
"00111111111111100000000000000011",	-- 1967: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 1968: 	addi	%sp, %sp, 4
"01011000000000000000010001010111",	-- 1969: 	jal	sin.2516
"10101011110111100000000000000100",	-- 1970: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 1971: 	lw	%ra, [%sp + 3]
"11001100000000010000000000000001",	-- 1972: 	lli	%r1, 1
"00111100001111100000000000000011",	-- 1973: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 1974: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 1975: 	addi	%sp, %sp, 5
"01011000000000000010101001001111",	-- 1976: 	jal	yj_fneg
"10101011110111100000000000000101",	-- 1977: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 1978: 	lw	%ra, [%sp + 4]
"00111011110000010000000000000011",	-- 1979: 	lw	%r1, [%sp + 3]
"00111011110000100000000000000001",	-- 1980: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 1981: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1982: 	sf	%f0, [%r1 + 0]
"00111111111111100000000000000100",	-- 1983: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 1984: 	addi	%sp, %sp, 5
"01011000000000000010101000111111",	-- 1985: 	jal	yj_read_float
"10101011110111100000000000000101",	-- 1986: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 1987: 	lw	%ra, [%sp + 4]
"00111111111111100000000000000100",	-- 1988: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 1989: 	addi	%sp, %sp, 5
"01011000000000000000011011000100",	-- 1990: 	jal	rad.2693
"10101011110111100000000000000101",	-- 1991: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 1992: 	lw	%ra, [%sp + 4]
"10010011110000010000000000000010",	-- 1993: 	lf	%f1, [%sp + 2]
"10110000000111100000000000000100",	-- 1994: 	sf	%f0, [%sp + 4]
"00001100001000000000000000000000",	-- 1995: 	movf	%f0, %f1
"00111111111111100000000000000101",	-- 1996: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 1997: 	addi	%sp, %sp, 6
"01011000000000000000010010010110",	-- 1998: 	jal	cos.2518
"10101011110111100000000000000110",	-- 1999: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 2000: 	lw	%ra, [%sp + 5]
"10010011110000010000000000000100",	-- 2001: 	lf	%f1, [%sp + 4]
"10110000000111100000000000000101",	-- 2002: 	sf	%f0, [%sp + 5]
"00001100001000000000000000000000",	-- 2003: 	movf	%f0, %f1
"00111111111111100000000000000110",	-- 2004: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 2005: 	addi	%sp, %sp, 7
"01011000000000000000010001010111",	-- 2006: 	jal	sin.2516
"10101011110111100000000000000111",	-- 2007: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 2008: 	lw	%ra, [%sp + 6]
"11001100000000010000000000000000",	-- 2009: 	lli	%r1, 0
"10010011110000010000000000000101",	-- 2010: 	lf	%f1, [%sp + 5]
"11101000001000000000000000000000",	-- 2011: 	mulf	%f0, %f1, %f0
"00111011110000100000000000000001",	-- 2012: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2013: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2014: 	sf	%f0, [%r1 + 0]
"10010011110000000000000000000100",	-- 2015: 	lf	%f0, [%sp + 4]
"00111111111111100000000000000110",	-- 2016: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 2017: 	addi	%sp, %sp, 7
"01011000000000000000010010010110",	-- 2018: 	jal	cos.2518
"10101011110111100000000000000111",	-- 2019: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 2020: 	lw	%ra, [%sp + 6]
"11001100000000010000000000000010",	-- 2021: 	lli	%r1, 2
"10010011110000010000000000000101",	-- 2022: 	lf	%f1, [%sp + 5]
"11101000001000000000000000000000",	-- 2023: 	mulf	%f0, %f1, %f0
"00111011110000100000000000000001",	-- 2024: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2025: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2026: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 2027: 	lli	%r1, 0
"00111100001111100000000000000110",	-- 2028: 	sw	%r1, [%sp + 6]
"00111111111111100000000000000111",	-- 2029: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 2030: 	addi	%sp, %sp, 8
"01011000000000000010101000111111",	-- 2031: 	jal	yj_read_float
"10101011110111100000000000001000",	-- 2032: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 2033: 	lw	%ra, [%sp + 7]
"00111011110000010000000000000110",	-- 2034: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000000",	-- 2035: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 2036: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2037: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 2038: 	jr	%ra
	-- rotate_quadratic_matrix.2699:
"11001100000000110000000000000000",	-- 2039: 	lli	%r3, 0
"10000100010000110001100000000000",	-- 2040: 	add	%r3, %r2, %r3
"10010000011000000000000000000000",	-- 2041: 	lf	%f0, [%r3 + 0]
"00111100001111100000000000000000",	-- 2042: 	sw	%r1, [%sp + 0]
"00111100010111100000000000000001",	-- 2043: 	sw	%r2, [%sp + 1]
"00111111111111100000000000000010",	-- 2044: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 2045: 	addi	%sp, %sp, 3
"01011000000000000000010010010110",	-- 2046: 	jal	cos.2518
"10101011110111100000000000000011",	-- 2047: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 2048: 	lw	%ra, [%sp + 2]
"11001100000000010000000000000000",	-- 2049: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 2050: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2051: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 2052: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000010",	-- 2053: 	sf	%f0, [%sp + 2]
"00001100001000000000000000000000",	-- 2054: 	movf	%f0, %f1
"00111111111111100000000000000011",	-- 2055: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 2056: 	addi	%sp, %sp, 4
"01011000000000000000010001010111",	-- 2057: 	jal	sin.2516
"10101011110111100000000000000100",	-- 2058: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 2059: 	lw	%ra, [%sp + 3]
"11001100000000010000000000000001",	-- 2060: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 2061: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2062: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 2063: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000011",	-- 2064: 	sf	%f0, [%sp + 3]
"00001100001000000000000000000000",	-- 2065: 	movf	%f0, %f1
"00111111111111100000000000000100",	-- 2066: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 2067: 	addi	%sp, %sp, 5
"01011000000000000000010010010110",	-- 2068: 	jal	cos.2518
"10101011110111100000000000000101",	-- 2069: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 2070: 	lw	%ra, [%sp + 4]
"11001100000000010000000000000001",	-- 2071: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 2072: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2073: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 2074: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000100",	-- 2075: 	sf	%f0, [%sp + 4]
"00001100001000000000000000000000",	-- 2076: 	movf	%f0, %f1
"00111111111111100000000000000101",	-- 2077: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 2078: 	addi	%sp, %sp, 6
"01011000000000000000010001010111",	-- 2079: 	jal	sin.2516
"10101011110111100000000000000110",	-- 2080: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 2081: 	lw	%ra, [%sp + 5]
"11001100000000010000000000000010",	-- 2082: 	lli	%r1, 2
"00111011110000100000000000000001",	-- 2083: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2084: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 2085: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000101",	-- 2086: 	sf	%f0, [%sp + 5]
"00001100001000000000000000000000",	-- 2087: 	movf	%f0, %f1
"00111111111111100000000000000110",	-- 2088: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 2089: 	addi	%sp, %sp, 7
"01011000000000000000010010010110",	-- 2090: 	jal	cos.2518
"10101011110111100000000000000111",	-- 2091: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 2092: 	lw	%ra, [%sp + 6]
"11001100000000010000000000000010",	-- 2093: 	lli	%r1, 2
"00111011110000100000000000000001",	-- 2094: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2095: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 2096: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000110",	-- 2097: 	sf	%f0, [%sp + 6]
"00001100001000000000000000000000",	-- 2098: 	movf	%f0, %f1
"00111111111111100000000000000111",	-- 2099: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 2100: 	addi	%sp, %sp, 8
"01011000000000000000010001010111",	-- 2101: 	jal	sin.2516
"10101011110111100000000000001000",	-- 2102: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 2103: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000110",	-- 2104: 	lf	%f1, [%sp + 6]
"10010011110000100000000000000100",	-- 2105: 	lf	%f2, [%sp + 4]
"11101000010000010001100000000000",	-- 2106: 	mulf	%f3, %f2, %f1
"10010011110001000000000000000101",	-- 2107: 	lf	%f4, [%sp + 5]
"10010011110001010000000000000011",	-- 2108: 	lf	%f5, [%sp + 3]
"11101000101001000011000000000000",	-- 2109: 	mulf	%f6, %f5, %f4
"11101000110000010011000000000000",	-- 2110: 	mulf	%f6, %f6, %f1
"10010011110001110000000000000010",	-- 2111: 	lf	%f7, [%sp + 2]
"11101000111000000100000000000000",	-- 2112: 	mulf	%f8, %f7, %f0
"11100100110010000011000000000000",	-- 2113: 	subf	%f6, %f6, %f8
"11101000111001000100000000000000",	-- 2114: 	mulf	%f8, %f7, %f4
"11101001000000010100000000000000",	-- 2115: 	mulf	%f8, %f8, %f1
"11101000101000000100100000000000",	-- 2116: 	mulf	%f9, %f5, %f0
"11100001000010010100000000000000",	-- 2117: 	addf	%f8, %f8, %f9
"11101000010000000100100000000000",	-- 2118: 	mulf	%f9, %f2, %f0
"11101000101001000101000000000000",	-- 2119: 	mulf	%f10, %f5, %f4
"11101001010000000101000000000000",	-- 2120: 	mulf	%f10, %f10, %f0
"11101000111000010101100000000000",	-- 2121: 	mulf	%f11, %f7, %f1
"11100001010010110101000000000000",	-- 2122: 	addf	%f10, %f10, %f11
"11101000111001000101100000000000",	-- 2123: 	mulf	%f11, %f7, %f4
"11101001011000000000000000000000",	-- 2124: 	mulf	%f0, %f11, %f0
"11101000101000010000100000000000",	-- 2125: 	mulf	%f1, %f5, %f1
"11100100000000010000000000000000",	-- 2126: 	subf	%f0, %f0, %f1
"10110000000111100000000000000111",	-- 2127: 	sf	%f0, [%sp + 7]
"10110001000111100000000000001000",	-- 2128: 	sf	%f8, [%sp + 8]
"10110001010111100000000000001001",	-- 2129: 	sf	%f10, [%sp + 9]
"10110000110111100000000000001010",	-- 2130: 	sf	%f6, [%sp + 10]
"10110001001111100000000000001011",	-- 2131: 	sf	%f9, [%sp + 11]
"10110000011111100000000000001100",	-- 2132: 	sf	%f3, [%sp + 12]
"00001100100000000000000000000000",	-- 2133: 	movf	%f0, %f4
"00111111111111100000000000001101",	-- 2134: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 2135: 	addi	%sp, %sp, 14
"01011000000000000010101001001111",	-- 2136: 	jal	yj_fneg
"10101011110111100000000000001110",	-- 2137: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 2138: 	lw	%ra, [%sp + 13]
"10010011110000010000000000000100",	-- 2139: 	lf	%f1, [%sp + 4]
"10010011110000100000000000000011",	-- 2140: 	lf	%f2, [%sp + 3]
"11101000010000010001000000000000",	-- 2141: 	mulf	%f2, %f2, %f1
"10010011110000110000000000000010",	-- 2142: 	lf	%f3, [%sp + 2]
"11101000011000010000100000000000",	-- 2143: 	mulf	%f1, %f3, %f1
"11001100000000010000000000000000",	-- 2144: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 2145: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 2146: 	add	%r1, %r2, %r1
"10010000001000110000000000000000",	-- 2147: 	lf	%f3, [%r1 + 0]
"11001100000000010000000000000001",	-- 2148: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 2149: 	add	%r1, %r2, %r1
"10010000001001000000000000000000",	-- 2150: 	lf	%f4, [%r1 + 0]
"11001100000000010000000000000010",	-- 2151: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 2152: 	add	%r1, %r2, %r1
"10010000001001010000000000000000",	-- 2153: 	lf	%f5, [%r1 + 0]
"11001100000000010000000000000000",	-- 2154: 	lli	%r1, 0
"10010011110001100000000000001100",	-- 2155: 	lf	%f6, [%sp + 12]
"10110000001111100000000000001101",	-- 2156: 	sf	%f1, [%sp + 13]
"10110000010111100000000000001110",	-- 2157: 	sf	%f2, [%sp + 14]
"00111100001111100000000000001111",	-- 2158: 	sw	%r1, [%sp + 15]
"10110000101111100000000000010000",	-- 2159: 	sf	%f5, [%sp + 16]
"10110000000111100000000000010001",	-- 2160: 	sf	%f0, [%sp + 17]
"10110000100111100000000000010010",	-- 2161: 	sf	%f4, [%sp + 18]
"10110000011111100000000000010011",	-- 2162: 	sf	%f3, [%sp + 19]
"00001100110000000000000000000000",	-- 2163: 	movf	%f0, %f6
"00111111111111100000000000010100",	-- 2164: 	sw	%ra, [%sp + 20]
"10100111110111100000000000010101",	-- 2165: 	addi	%sp, %sp, 21
"01011000000000000000010011101111",	-- 2166: 	jal	fsqr.2530
"10101011110111100000000000010101",	-- 2167: 	subi	%sp, %sp, 21
"00111011110111110000000000010100",	-- 2168: 	lw	%ra, [%sp + 20]
"10010011110000010000000000010011",	-- 2169: 	lf	%f1, [%sp + 19]
"11101000001000000000000000000000",	-- 2170: 	mulf	%f0, %f1, %f0
"10010011110000100000000000001011",	-- 2171: 	lf	%f2, [%sp + 11]
"10110000000111100000000000010100",	-- 2172: 	sf	%f0, [%sp + 20]
"00001100010000000000000000000000",	-- 2173: 	movf	%f0, %f2
"00111111111111100000000000010101",	-- 2174: 	sw	%ra, [%sp + 21]
"10100111110111100000000000010110",	-- 2175: 	addi	%sp, %sp, 22
"01011000000000000000010011101111",	-- 2176: 	jal	fsqr.2530
"10101011110111100000000000010110",	-- 2177: 	subi	%sp, %sp, 22
"00111011110111110000000000010101",	-- 2178: 	lw	%ra, [%sp + 21]
"10010011110000010000000000010010",	-- 2179: 	lf	%f1, [%sp + 18]
"11101000001000000000000000000000",	-- 2180: 	mulf	%f0, %f1, %f0
"10010011110000100000000000010100",	-- 2181: 	lf	%f2, [%sp + 20]
"11100000010000000000000000000000",	-- 2182: 	addf	%f0, %f2, %f0
"10010011110000100000000000010001",	-- 2183: 	lf	%f2, [%sp + 17]
"10110000000111100000000000010101",	-- 2184: 	sf	%f0, [%sp + 21]
"00001100010000000000000000000000",	-- 2185: 	movf	%f0, %f2
"00111111111111100000000000010110",	-- 2186: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 2187: 	addi	%sp, %sp, 23
"01011000000000000000010011101111",	-- 2188: 	jal	fsqr.2530
"10101011110111100000000000010111",	-- 2189: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 2190: 	lw	%ra, [%sp + 22]
"10010011110000010000000000010000",	-- 2191: 	lf	%f1, [%sp + 16]
"11101000001000000000000000000000",	-- 2192: 	mulf	%f0, %f1, %f0
"10010011110000100000000000010101",	-- 2193: 	lf	%f2, [%sp + 21]
"11100000010000000000000000000000",	-- 2194: 	addf	%f0, %f2, %f0
"00111011110000010000000000001111",	-- 2195: 	lw	%r1, [%sp + 15]
"00111011110000100000000000000000",	-- 2196: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 2197: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2198: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2199: 	lli	%r1, 1
"10010011110000000000000000001010",	-- 2200: 	lf	%f0, [%sp + 10]
"00111100001111100000000000010110",	-- 2201: 	sw	%r1, [%sp + 22]
"00111111111111100000000000010111",	-- 2202: 	sw	%ra, [%sp + 23]
"10100111110111100000000000011000",	-- 2203: 	addi	%sp, %sp, 24
"01011000000000000000010011101111",	-- 2204: 	jal	fsqr.2530
"10101011110111100000000000011000",	-- 2205: 	subi	%sp, %sp, 24
"00111011110111110000000000010111",	-- 2206: 	lw	%ra, [%sp + 23]
"10010011110000010000000000010011",	-- 2207: 	lf	%f1, [%sp + 19]
"11101000001000000000000000000000",	-- 2208: 	mulf	%f0, %f1, %f0
"10010011110000100000000000001001",	-- 2209: 	lf	%f2, [%sp + 9]
"10110000000111100000000000010111",	-- 2210: 	sf	%f0, [%sp + 23]
"00001100010000000000000000000000",	-- 2211: 	movf	%f0, %f2
"00111111111111100000000000011000",	-- 2212: 	sw	%ra, [%sp + 24]
"10100111110111100000000000011001",	-- 2213: 	addi	%sp, %sp, 25
"01011000000000000000010011101111",	-- 2214: 	jal	fsqr.2530
"10101011110111100000000000011001",	-- 2215: 	subi	%sp, %sp, 25
"00111011110111110000000000011000",	-- 2216: 	lw	%ra, [%sp + 24]
"10010011110000010000000000010010",	-- 2217: 	lf	%f1, [%sp + 18]
"11101000001000000000000000000000",	-- 2218: 	mulf	%f0, %f1, %f0
"10010011110000100000000000010111",	-- 2219: 	lf	%f2, [%sp + 23]
"11100000010000000000000000000000",	-- 2220: 	addf	%f0, %f2, %f0
"10010011110000100000000000001110",	-- 2221: 	lf	%f2, [%sp + 14]
"10110000000111100000000000011000",	-- 2222: 	sf	%f0, [%sp + 24]
"00001100010000000000000000000000",	-- 2223: 	movf	%f0, %f2
"00111111111111100000000000011001",	-- 2224: 	sw	%ra, [%sp + 25]
"10100111110111100000000000011010",	-- 2225: 	addi	%sp, %sp, 26
"01011000000000000000010011101111",	-- 2226: 	jal	fsqr.2530
"10101011110111100000000000011010",	-- 2227: 	subi	%sp, %sp, 26
"00111011110111110000000000011001",	-- 2228: 	lw	%ra, [%sp + 25]
"10010011110000010000000000010000",	-- 2229: 	lf	%f1, [%sp + 16]
"11101000001000000000000000000000",	-- 2230: 	mulf	%f0, %f1, %f0
"10010011110000100000000000011000",	-- 2231: 	lf	%f2, [%sp + 24]
"11100000010000000000000000000000",	-- 2232: 	addf	%f0, %f2, %f0
"00111011110000010000000000010110",	-- 2233: 	lw	%r1, [%sp + 22]
"00111011110000100000000000000000",	-- 2234: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 2235: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2236: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2237: 	lli	%r1, 2
"10010011110000000000000000001000",	-- 2238: 	lf	%f0, [%sp + 8]
"00111100001111100000000000011001",	-- 2239: 	sw	%r1, [%sp + 25]
"00111111111111100000000000011010",	-- 2240: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 2241: 	addi	%sp, %sp, 27
"01011000000000000000010011101111",	-- 2242: 	jal	fsqr.2530
"10101011110111100000000000011011",	-- 2243: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 2244: 	lw	%ra, [%sp + 26]
"10010011110000010000000000010011",	-- 2245: 	lf	%f1, [%sp + 19]
"11101000001000000000000000000000",	-- 2246: 	mulf	%f0, %f1, %f0
"10010011110000100000000000000111",	-- 2247: 	lf	%f2, [%sp + 7]
"10110000000111100000000000011010",	-- 2248: 	sf	%f0, [%sp + 26]
"00001100010000000000000000000000",	-- 2249: 	movf	%f0, %f2
"00111111111111100000000000011011",	-- 2250: 	sw	%ra, [%sp + 27]
"10100111110111100000000000011100",	-- 2251: 	addi	%sp, %sp, 28
"01011000000000000000010011101111",	-- 2252: 	jal	fsqr.2530
"10101011110111100000000000011100",	-- 2253: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 2254: 	lw	%ra, [%sp + 27]
"10010011110000010000000000010010",	-- 2255: 	lf	%f1, [%sp + 18]
"11101000001000000000000000000000",	-- 2256: 	mulf	%f0, %f1, %f0
"10010011110000100000000000011010",	-- 2257: 	lf	%f2, [%sp + 26]
"11100000010000000000000000000000",	-- 2258: 	addf	%f0, %f2, %f0
"10010011110000100000000000001101",	-- 2259: 	lf	%f2, [%sp + 13]
"10110000000111100000000000011011",	-- 2260: 	sf	%f0, [%sp + 27]
"00001100010000000000000000000000",	-- 2261: 	movf	%f0, %f2
"00111111111111100000000000011100",	-- 2262: 	sw	%ra, [%sp + 28]
"10100111110111100000000000011101",	-- 2263: 	addi	%sp, %sp, 29
"01011000000000000000010011101111",	-- 2264: 	jal	fsqr.2530
"10101011110111100000000000011101",	-- 2265: 	subi	%sp, %sp, 29
"00111011110111110000000000011100",	-- 2266: 	lw	%ra, [%sp + 28]
"10010011110000010000000000010000",	-- 2267: 	lf	%f1, [%sp + 16]
"11101000001000000000000000000000",	-- 2268: 	mulf	%f0, %f1, %f0
"10010011110000100000000000011011",	-- 2269: 	lf	%f2, [%sp + 27]
"11100000010000000000000000000000",	-- 2270: 	addf	%f0, %f2, %f0
"00111011110000010000000000011001",	-- 2271: 	lw	%r1, [%sp + 25]
"00111011110000100000000000000000",	-- 2272: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 2273: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2274: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 2275: 	lli	%r1, 0
"00010100000000000000000000000000",	-- 2276: 	llif	%f0, 2.000000
"00010000000000000100000000000000",	-- 2277: 	lhif	%f0, 2.000000
"10010011110000100000000000001010",	-- 2278: 	lf	%f2, [%sp + 10]
"10010011110000110000000000010011",	-- 2279: 	lf	%f3, [%sp + 19]
"11101000011000100010000000000000",	-- 2280: 	mulf	%f4, %f3, %f2
"10010011110001010000000000001000",	-- 2281: 	lf	%f5, [%sp + 8]
"11101000100001010010000000000000",	-- 2282: 	mulf	%f4, %f4, %f5
"10010011110001100000000000001001",	-- 2283: 	lf	%f6, [%sp + 9]
"10010011110001110000000000010010",	-- 2284: 	lf	%f7, [%sp + 18]
"11101000111001100100000000000000",	-- 2285: 	mulf	%f8, %f7, %f6
"10010011110010010000000000000111",	-- 2286: 	lf	%f9, [%sp + 7]
"11101001000010010100000000000000",	-- 2287: 	mulf	%f8, %f8, %f9
"11100000100010000010000000000000",	-- 2288: 	addf	%f4, %f4, %f8
"10010011110010000000000000001110",	-- 2289: 	lf	%f8, [%sp + 14]
"11101000001010000101000000000000",	-- 2290: 	mulf	%f10, %f1, %f8
"10010011110010110000000000001101",	-- 2291: 	lf	%f11, [%sp + 13]
"11101001010010110101000000000000",	-- 2292: 	mulf	%f10, %f10, %f11
"11100000100010100010000000000000",	-- 2293: 	addf	%f4, %f4, %f10
"11101000000001000000000000000000",	-- 2294: 	mulf	%f0, %f0, %f4
"00111011110000100000000000000001",	-- 2295: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2296: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2297: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2298: 	lli	%r1, 1
"00010100000000000000000000000000",	-- 2299: 	llif	%f0, 2.000000
"00010000000000000100000000000000",	-- 2300: 	lhif	%f0, 2.000000
"10010011110001000000000000001100",	-- 2301: 	lf	%f4, [%sp + 12]
"11101000011001000101000000000000",	-- 2302: 	mulf	%f10, %f3, %f4
"11101001010001010010100000000000",	-- 2303: 	mulf	%f5, %f10, %f5
"10010011110010100000000000001011",	-- 2304: 	lf	%f10, [%sp + 11]
"11101000111010100110000000000000",	-- 2305: 	mulf	%f12, %f7, %f10
"11101001100010010100100000000000",	-- 2306: 	mulf	%f9, %f12, %f9
"11100000101010010010100000000000",	-- 2307: 	addf	%f5, %f5, %f9
"10010011110010010000000000010001",	-- 2308: 	lf	%f9, [%sp + 17]
"11101000001010010110000000000000",	-- 2309: 	mulf	%f12, %f1, %f9
"11101001100010110101100000000000",	-- 2310: 	mulf	%f11, %f12, %f11
"11100000101010110010100000000000",	-- 2311: 	addf	%f5, %f5, %f11
"11101000000001010000000000000000",	-- 2312: 	mulf	%f0, %f0, %f5
"10000100010000010000100000000000",	-- 2313: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2314: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2315: 	lli	%r1, 2
"00010100000000000000000000000000",	-- 2316: 	llif	%f0, 2.000000
"00010000000000000100000000000000",	-- 2317: 	lhif	%f0, 2.000000
"11101000011001000001100000000000",	-- 2318: 	mulf	%f3, %f3, %f4
"11101000011000100001000000000000",	-- 2319: 	mulf	%f2, %f3, %f2
"11101000111010100001100000000000",	-- 2320: 	mulf	%f3, %f7, %f10
"11101000011001100001100000000000",	-- 2321: 	mulf	%f3, %f3, %f6
"11100000010000110001000000000000",	-- 2322: 	addf	%f2, %f2, %f3
"11101000001010010000100000000000",	-- 2323: 	mulf	%f1, %f1, %f9
"11101000001010000000100000000000",	-- 2324: 	mulf	%f1, %f1, %f8
"11100000010000010000100000000000",	-- 2325: 	addf	%f1, %f2, %f1
"11101000000000010000000000000000",	-- 2326: 	mulf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 2327: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2328: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 2329: 	jr	%ra
	-- read_nth_object.2702:
"00111011011000100000000000000001",	-- 2330: 	lw	%r2, [%r27 + 1]
"00111100001111100000000000000000",	-- 2331: 	sw	%r1, [%sp + 0]
"00111100010111100000000000000001",	-- 2332: 	sw	%r2, [%sp + 1]
"00111111111111100000000000000010",	-- 2333: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 2334: 	addi	%sp, %sp, 3
"01011000000000000010101000110010",	-- 2335: 	jal	yj_read_int
"10101011110111100000000000000011",	-- 2336: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 2337: 	lw	%ra, [%sp + 2]
"11001100000000101111111111111111",	-- 2338: 	lli	%r2, -1
"11001000000000101111111111111111",	-- 2339: 	lhi	%r2, -1
"00101000001000100000000000000011",	-- 2340: 	bneq	%r1, %r2, bneq_else.8961
"11001100000000010000000000000000",	-- 2341: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 2342: 	jr	%ra
	-- bneq_else.8961:
"00111100001111100000000000000010",	-- 2343: 	sw	%r1, [%sp + 2]
"00111111111111100000000000000011",	-- 2344: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 2345: 	addi	%sp, %sp, 4
"01011000000000000010101000110010",	-- 2346: 	jal	yj_read_int
"10101011110111100000000000000100",	-- 2347: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 2348: 	lw	%ra, [%sp + 3]
"00111100001111100000000000000011",	-- 2349: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 2350: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 2351: 	addi	%sp, %sp, 5
"01011000000000000010101000110010",	-- 2352: 	jal	yj_read_int
"10101011110111100000000000000101",	-- 2353: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 2354: 	lw	%ra, [%sp + 4]
"00111100001111100000000000000100",	-- 2355: 	sw	%r1, [%sp + 4]
"00111111111111100000000000000101",	-- 2356: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 2357: 	addi	%sp, %sp, 6
"01011000000000000010101000110010",	-- 2358: 	jal	yj_read_int
"10101011110111100000000000000110",	-- 2359: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 2360: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000011",	-- 2361: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 2362: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2363: 	lhif	%f0, 0.000000
"00111100001111100000000000000101",	-- 2364: 	sw	%r1, [%sp + 5]
"10000100000000100000100000000000",	-- 2365: 	add	%r1, %r0, %r2
"00111111111111100000000000000110",	-- 2366: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 2367: 	addi	%sp, %sp, 7
"01011000000000000010101000100010",	-- 2368: 	jal	yj_create_float_array
"10101011110111100000000000000111",	-- 2369: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 2370: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 2371: 	lli	%r2, 0
"00111100010111100000000000000110",	-- 2372: 	sw	%r2, [%sp + 6]
"00111100001111100000000000000111",	-- 2373: 	sw	%r1, [%sp + 7]
"00111111111111100000000000001000",	-- 2374: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 2375: 	addi	%sp, %sp, 9
"01011000000000000010101000111111",	-- 2376: 	jal	yj_read_float
"10101011110111100000000000001001",	-- 2377: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 2378: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000110",	-- 2379: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000111",	-- 2380: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 2381: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2382: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2383: 	lli	%r1, 1
"00111100001111100000000000001000",	-- 2384: 	sw	%r1, [%sp + 8]
"00111111111111100000000000001001",	-- 2385: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 2386: 	addi	%sp, %sp, 10
"01011000000000000010101000111111",	-- 2387: 	jal	yj_read_float
"10101011110111100000000000001010",	-- 2388: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 2389: 	lw	%ra, [%sp + 9]
"00111011110000010000000000001000",	-- 2390: 	lw	%r1, [%sp + 8]
"00111011110000100000000000000111",	-- 2391: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 2392: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2393: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2394: 	lli	%r1, 2
"00111100001111100000000000001001",	-- 2395: 	sw	%r1, [%sp + 9]
"00111111111111100000000000001010",	-- 2396: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 2397: 	addi	%sp, %sp, 11
"01011000000000000010101000111111",	-- 2398: 	jal	yj_read_float
"10101011110111100000000000001011",	-- 2399: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 2400: 	lw	%ra, [%sp + 10]
"00111011110000010000000000001001",	-- 2401: 	lw	%r1, [%sp + 9]
"00111011110000100000000000000111",	-- 2402: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 2403: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2404: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 2405: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 2406: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2407: 	lhif	%f0, 0.000000
"00111111111111100000000000001010",	-- 2408: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 2409: 	addi	%sp, %sp, 11
"01011000000000000010101000100010",	-- 2410: 	jal	yj_create_float_array
"10101011110111100000000000001011",	-- 2411: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 2412: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 2413: 	lli	%r2, 0
"00111100010111100000000000001010",	-- 2414: 	sw	%r2, [%sp + 10]
"00111100001111100000000000001011",	-- 2415: 	sw	%r1, [%sp + 11]
"00111111111111100000000000001100",	-- 2416: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 2417: 	addi	%sp, %sp, 13
"01011000000000000010101000111111",	-- 2418: 	jal	yj_read_float
"10101011110111100000000000001101",	-- 2419: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 2420: 	lw	%ra, [%sp + 12]
"00111011110000010000000000001010",	-- 2421: 	lw	%r1, [%sp + 10]
"00111011110000100000000000001011",	-- 2422: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 2423: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2424: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2425: 	lli	%r1, 1
"00111100001111100000000000001100",	-- 2426: 	sw	%r1, [%sp + 12]
"00111111111111100000000000001101",	-- 2427: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 2428: 	addi	%sp, %sp, 14
"01011000000000000010101000111111",	-- 2429: 	jal	yj_read_float
"10101011110111100000000000001110",	-- 2430: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 2431: 	lw	%ra, [%sp + 13]
"00111011110000010000000000001100",	-- 2432: 	lw	%r1, [%sp + 12]
"00111011110000100000000000001011",	-- 2433: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 2434: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2435: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2436: 	lli	%r1, 2
"00111100001111100000000000001101",	-- 2437: 	sw	%r1, [%sp + 13]
"00111111111111100000000000001110",	-- 2438: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 2439: 	addi	%sp, %sp, 15
"01011000000000000010101000111111",	-- 2440: 	jal	yj_read_float
"10101011110111100000000000001111",	-- 2441: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 2442: 	lw	%ra, [%sp + 14]
"00111011110000010000000000001101",	-- 2443: 	lw	%r1, [%sp + 13]
"00111011110000100000000000001011",	-- 2444: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 2445: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2446: 	sf	%f0, [%r1 + 0]
"00111111111111100000000000001110",	-- 2447: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 2448: 	addi	%sp, %sp, 15
"01011000000000000010101000111111",	-- 2449: 	jal	yj_read_float
"10101011110111100000000000001111",	-- 2450: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 2451: 	lw	%ra, [%sp + 14]
"00111111111111100000000000001110",	-- 2452: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 2453: 	addi	%sp, %sp, 15
"01011000000000000000010011011011",	-- 2454: 	jal	fisneg.2524
"10101011110111100000000000001111",	-- 2455: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 2456: 	lw	%ra, [%sp + 14]
"11001100000000100000000000000010",	-- 2457: 	lli	%r2, 2
"00010100000000000000000000000000",	-- 2458: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2459: 	lhif	%f0, 0.000000
"00111100001111100000000000001110",	-- 2460: 	sw	%r1, [%sp + 14]
"10000100000000100000100000000000",	-- 2461: 	add	%r1, %r0, %r2
"00111111111111100000000000001111",	-- 2462: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 2463: 	addi	%sp, %sp, 16
"01011000000000000010101000100010",	-- 2464: 	jal	yj_create_float_array
"10101011110111100000000000010000",	-- 2465: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 2466: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 2467: 	lli	%r2, 0
"00111100010111100000000000001111",	-- 2468: 	sw	%r2, [%sp + 15]
"00111100001111100000000000010000",	-- 2469: 	sw	%r1, [%sp + 16]
"00111111111111100000000000010001",	-- 2470: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 2471: 	addi	%sp, %sp, 18
"01011000000000000010101000111111",	-- 2472: 	jal	yj_read_float
"10101011110111100000000000010010",	-- 2473: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 2474: 	lw	%ra, [%sp + 17]
"00111011110000010000000000001111",	-- 2475: 	lw	%r1, [%sp + 15]
"00111011110000100000000000010000",	-- 2476: 	lw	%r2, [%sp + 16]
"10000100010000010000100000000000",	-- 2477: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2478: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2479: 	lli	%r1, 1
"00111100001111100000000000010001",	-- 2480: 	sw	%r1, [%sp + 17]
"00111111111111100000000000010010",	-- 2481: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 2482: 	addi	%sp, %sp, 19
"01011000000000000010101000111111",	-- 2483: 	jal	yj_read_float
"10101011110111100000000000010011",	-- 2484: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 2485: 	lw	%ra, [%sp + 18]
"00111011110000010000000000010001",	-- 2486: 	lw	%r1, [%sp + 17]
"00111011110000100000000000010000",	-- 2487: 	lw	%r2, [%sp + 16]
"10000100010000010000100000000000",	-- 2488: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2489: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 2490: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 2491: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2492: 	lhif	%f0, 0.000000
"00111111111111100000000000010010",	-- 2493: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 2494: 	addi	%sp, %sp, 19
"01011000000000000010101000100010",	-- 2495: 	jal	yj_create_float_array
"10101011110111100000000000010011",	-- 2496: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 2497: 	lw	%ra, [%sp + 18]
"11001100000000100000000000000000",	-- 2498: 	lli	%r2, 0
"00111100010111100000000000010010",	-- 2499: 	sw	%r2, [%sp + 18]
"00111100001111100000000000010011",	-- 2500: 	sw	%r1, [%sp + 19]
"00111111111111100000000000010100",	-- 2501: 	sw	%ra, [%sp + 20]
"10100111110111100000000000010101",	-- 2502: 	addi	%sp, %sp, 21
"01011000000000000010101000111111",	-- 2503: 	jal	yj_read_float
"10101011110111100000000000010101",	-- 2504: 	subi	%sp, %sp, 21
"00111011110111110000000000010100",	-- 2505: 	lw	%ra, [%sp + 20]
"00111011110000010000000000010010",	-- 2506: 	lw	%r1, [%sp + 18]
"00111011110000100000000000010011",	-- 2507: 	lw	%r2, [%sp + 19]
"10000100010000010000100000000000",	-- 2508: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2509: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2510: 	lli	%r1, 1
"00111100001111100000000000010100",	-- 2511: 	sw	%r1, [%sp + 20]
"00111111111111100000000000010101",	-- 2512: 	sw	%ra, [%sp + 21]
"10100111110111100000000000010110",	-- 2513: 	addi	%sp, %sp, 22
"01011000000000000010101000111111",	-- 2514: 	jal	yj_read_float
"10101011110111100000000000010110",	-- 2515: 	subi	%sp, %sp, 22
"00111011110111110000000000010101",	-- 2516: 	lw	%ra, [%sp + 21]
"00111011110000010000000000010100",	-- 2517: 	lw	%r1, [%sp + 20]
"00111011110000100000000000010011",	-- 2518: 	lw	%r2, [%sp + 19]
"10000100010000010000100000000000",	-- 2519: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2520: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2521: 	lli	%r1, 2
"00111100001111100000000000010101",	-- 2522: 	sw	%r1, [%sp + 21]
"00111111111111100000000000010110",	-- 2523: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 2524: 	addi	%sp, %sp, 23
"01011000000000000010101000111111",	-- 2525: 	jal	yj_read_float
"10101011110111100000000000010111",	-- 2526: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 2527: 	lw	%ra, [%sp + 22]
"00111011110000010000000000010101",	-- 2528: 	lw	%r1, [%sp + 21]
"00111011110000100000000000010011",	-- 2529: 	lw	%r2, [%sp + 19]
"10000100010000010000100000000000",	-- 2530: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2531: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 2532: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 2533: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2534: 	lhif	%f0, 0.000000
"00111111111111100000000000010110",	-- 2535: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 2536: 	addi	%sp, %sp, 23
"01011000000000000010101000100010",	-- 2537: 	jal	yj_create_float_array
"10101011110111100000000000010111",	-- 2538: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 2539: 	lw	%ra, [%sp + 22]
"11001100000000100000000000000000",	-- 2540: 	lli	%r2, 0
"00111011110000110000000000000101",	-- 2541: 	lw	%r3, [%sp + 5]
"00111100001111100000000000010110",	-- 2542: 	sw	%r1, [%sp + 22]
"00101000011000100000000000000010",	-- 2543: 	bneq	%r3, %r2, bneq_else.8962
"01010100000000000000101000100001",	-- 2544: 	j	bneq_cont.8963
	-- bneq_else.8962:
"11001100000000100000000000000000",	-- 2545: 	lli	%r2, 0
"00111100010111100000000000010111",	-- 2546: 	sw	%r2, [%sp + 23]
"00111111111111100000000000011000",	-- 2547: 	sw	%ra, [%sp + 24]
"10100111110111100000000000011001",	-- 2548: 	addi	%sp, %sp, 25
"01011000000000000010101000111111",	-- 2549: 	jal	yj_read_float
"10101011110111100000000000011001",	-- 2550: 	subi	%sp, %sp, 25
"00111011110111110000000000011000",	-- 2551: 	lw	%ra, [%sp + 24]
"00111111111111100000000000011000",	-- 2552: 	sw	%ra, [%sp + 24]
"10100111110111100000000000011001",	-- 2553: 	addi	%sp, %sp, 25
"01011000000000000000011011000100",	-- 2554: 	jal	rad.2693
"10101011110111100000000000011001",	-- 2555: 	subi	%sp, %sp, 25
"00111011110111110000000000011000",	-- 2556: 	lw	%ra, [%sp + 24]
"00111011110000010000000000010111",	-- 2557: 	lw	%r1, [%sp + 23]
"00111011110000100000000000010110",	-- 2558: 	lw	%r2, [%sp + 22]
"10000100010000010000100000000000",	-- 2559: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2560: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2561: 	lli	%r1, 1
"00111100001111100000000000011000",	-- 2562: 	sw	%r1, [%sp + 24]
"00111111111111100000000000011001",	-- 2563: 	sw	%ra, [%sp + 25]
"10100111110111100000000000011010",	-- 2564: 	addi	%sp, %sp, 26
"01011000000000000010101000111111",	-- 2565: 	jal	yj_read_float
"10101011110111100000000000011010",	-- 2566: 	subi	%sp, %sp, 26
"00111011110111110000000000011001",	-- 2567: 	lw	%ra, [%sp + 25]
"00111111111111100000000000011001",	-- 2568: 	sw	%ra, [%sp + 25]
"10100111110111100000000000011010",	-- 2569: 	addi	%sp, %sp, 26
"01011000000000000000011011000100",	-- 2570: 	jal	rad.2693
"10101011110111100000000000011010",	-- 2571: 	subi	%sp, %sp, 26
"00111011110111110000000000011001",	-- 2572: 	lw	%ra, [%sp + 25]
"00111011110000010000000000011000",	-- 2573: 	lw	%r1, [%sp + 24]
"00111011110000100000000000010110",	-- 2574: 	lw	%r2, [%sp + 22]
"10000100010000010000100000000000",	-- 2575: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2576: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2577: 	lli	%r1, 2
"00111100001111100000000000011001",	-- 2578: 	sw	%r1, [%sp + 25]
"00111111111111100000000000011010",	-- 2579: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 2580: 	addi	%sp, %sp, 27
"01011000000000000010101000111111",	-- 2581: 	jal	yj_read_float
"10101011110111100000000000011011",	-- 2582: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 2583: 	lw	%ra, [%sp + 26]
"00111111111111100000000000011010",	-- 2584: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 2585: 	addi	%sp, %sp, 27
"01011000000000000000011011000100",	-- 2586: 	jal	rad.2693
"10101011110111100000000000011011",	-- 2587: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 2588: 	lw	%ra, [%sp + 26]
"00111011110000010000000000011001",	-- 2589: 	lw	%r1, [%sp + 25]
"00111011110000100000000000010110",	-- 2590: 	lw	%r2, [%sp + 22]
"10000100010000010000100000000000",	-- 2591: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2592: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.8963:
"11001100000000010000000000000010",	-- 2593: 	lli	%r1, 2
"00111011110000100000000000000011",	-- 2594: 	lw	%r2, [%sp + 3]
"00101000010000010000000000000011",	-- 2595: 	bneq	%r2, %r1, bneq_else.8964
"11001100000000010000000000000001",	-- 2596: 	lli	%r1, 1
"01010100000000000000101000100111",	-- 2597: 	j	bneq_cont.8965
	-- bneq_else.8964:
"00111011110000010000000000001110",	-- 2598: 	lw	%r1, [%sp + 14]
	-- bneq_cont.8965:
"11001100000000110000000000000100",	-- 2599: 	lli	%r3, 4
"00010100000000000000000000000000",	-- 2600: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2601: 	lhif	%f0, 0.000000
"00111100001111100000000000011010",	-- 2602: 	sw	%r1, [%sp + 26]
"10000100000000110000100000000000",	-- 2603: 	add	%r1, %r0, %r3
"00111111111111100000000000011011",	-- 2604: 	sw	%ra, [%sp + 27]
"10100111110111100000000000011100",	-- 2605: 	addi	%sp, %sp, 28
"01011000000000000010101000100010",	-- 2606: 	jal	yj_create_float_array
"10101011110111100000000000011100",	-- 2607: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 2608: 	lw	%ra, [%sp + 27]
"10000100000111010001000000000000",	-- 2609: 	add	%r2, %r0, %hp
"10100111101111010000000000001011",	-- 2610: 	addi	%hp, %hp, 11
"00111100001000100000000000001010",	-- 2611: 	sw	%r1, [%r2 + 10]
"00111011110000010000000000010110",	-- 2612: 	lw	%r1, [%sp + 22]
"00111100001000100000000000001001",	-- 2613: 	sw	%r1, [%r2 + 9]
"00111011110000110000000000010011",	-- 2614: 	lw	%r3, [%sp + 19]
"00111100011000100000000000001000",	-- 2615: 	sw	%r3, [%r2 + 8]
"00111011110000110000000000010000",	-- 2616: 	lw	%r3, [%sp + 16]
"00111100011000100000000000000111",	-- 2617: 	sw	%r3, [%r2 + 7]
"00111011110000110000000000011010",	-- 2618: 	lw	%r3, [%sp + 26]
"00111100011000100000000000000110",	-- 2619: 	sw	%r3, [%r2 + 6]
"00111011110000110000000000001011",	-- 2620: 	lw	%r3, [%sp + 11]
"00111100011000100000000000000101",	-- 2621: 	sw	%r3, [%r2 + 5]
"00111011110000110000000000000111",	-- 2622: 	lw	%r3, [%sp + 7]
"00111100011000100000000000000100",	-- 2623: 	sw	%r3, [%r2 + 4]
"00111011110001000000000000000101",	-- 2624: 	lw	%r4, [%sp + 5]
"00111100100000100000000000000011",	-- 2625: 	sw	%r4, [%r2 + 3]
"00111011110001010000000000000100",	-- 2626: 	lw	%r5, [%sp + 4]
"00111100101000100000000000000010",	-- 2627: 	sw	%r5, [%r2 + 2]
"00111011110001010000000000000011",	-- 2628: 	lw	%r5, [%sp + 3]
"00111100101000100000000000000001",	-- 2629: 	sw	%r5, [%r2 + 1]
"00111011110001100000000000000010",	-- 2630: 	lw	%r6, [%sp + 2]
"00111100110000100000000000000000",	-- 2631: 	sw	%r6, [%r2 + 0]
"00111011110001100000000000000000",	-- 2632: 	lw	%r6, [%sp + 0]
"00111011110001110000000000000001",	-- 2633: 	lw	%r7, [%sp + 1]
"10000100111001100011000000000000",	-- 2634: 	add	%r6, %r7, %r6
"00111100010001100000000000000000",	-- 2635: 	sw	%r2, [%r6 + 0]
"11001100000000100000000000000011",	-- 2636: 	lli	%r2, 3
"00101000101000100000000001101110",	-- 2637: 	bneq	%r5, %r2, bneq_else.8966
"11001100000000100000000000000000",	-- 2638: 	lli	%r2, 0
"10000100011000100001000000000000",	-- 2639: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 2640: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000000",	-- 2641: 	lli	%r2, 0
"00111100010111100000000000011011",	-- 2642: 	sw	%r2, [%sp + 27]
"10110000000111100000000000011100",	-- 2643: 	sf	%f0, [%sp + 28]
"00111111111111100000000000011101",	-- 2644: 	sw	%ra, [%sp + 29]
"10100111110111100000000000011110",	-- 2645: 	addi	%sp, %sp, 30
"01011000000000000000010011100010",	-- 2646: 	jal	fiszero.2526
"10101011110111100000000000011110",	-- 2647: 	subi	%sp, %sp, 30
"00111011110111110000000000011101",	-- 2648: 	lw	%ra, [%sp + 29]
"11001100000000100000000000000000",	-- 2649: 	lli	%r2, 0
"00101000001000100000000000010010",	-- 2650: 	bneq	%r1, %r2, bneq_else.8968
"10010011110000000000000000011100",	-- 2651: 	lf	%f0, [%sp + 28]
"00111111111111100000000000011101",	-- 2652: 	sw	%ra, [%sp + 29]
"10100111110111100000000000011110",	-- 2653: 	addi	%sp, %sp, 30
"01011000000000000000010100000000",	-- 2654: 	jal	sgn.2568
"10101011110111100000000000011110",	-- 2655: 	subi	%sp, %sp, 30
"00111011110111110000000000011101",	-- 2656: 	lw	%ra, [%sp + 29]
"10010011110000010000000000011100",	-- 2657: 	lf	%f1, [%sp + 28]
"10110000000111100000000000011101",	-- 2658: 	sf	%f0, [%sp + 29]
"00001100001000000000000000000000",	-- 2659: 	movf	%f0, %f1
"00111111111111100000000000011110",	-- 2660: 	sw	%ra, [%sp + 30]
"10100111110111100000000000011111",	-- 2661: 	addi	%sp, %sp, 31
"01011000000000000000010011101111",	-- 2662: 	jal	fsqr.2530
"10101011110111100000000000011111",	-- 2663: 	subi	%sp, %sp, 31
"00111011110111110000000000011110",	-- 2664: 	lw	%ra, [%sp + 30]
"10010011110000010000000000011101",	-- 2665: 	lf	%f1, [%sp + 29]
"11101100001000000000000000000000",	-- 2666: 	divf	%f0, %f1, %f0
"01010100000000000000101001101110",	-- 2667: 	j	bneq_cont.8969
	-- bneq_else.8968:
"00010100000000000000000000000000",	-- 2668: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2669: 	lhif	%f0, 0.000000
	-- bneq_cont.8969:
"00111011110000010000000000011011",	-- 2670: 	lw	%r1, [%sp + 27]
"00111011110000100000000000000111",	-- 2671: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 2672: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2673: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2674: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 2675: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 2676: 	lf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2677: 	lli	%r1, 1
"00111100001111100000000000011110",	-- 2678: 	sw	%r1, [%sp + 30]
"10110000000111100000000000011111",	-- 2679: 	sf	%f0, [%sp + 31]
"00111111111111100000000000100000",	-- 2680: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 2681: 	addi	%sp, %sp, 33
"01011000000000000000010011100010",	-- 2682: 	jal	fiszero.2526
"10101011110111100000000000100001",	-- 2683: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 2684: 	lw	%ra, [%sp + 32]
"11001100000000100000000000000000",	-- 2685: 	lli	%r2, 0
"00101000001000100000000000010010",	-- 2686: 	bneq	%r1, %r2, bneq_else.8970
"10010011110000000000000000011111",	-- 2687: 	lf	%f0, [%sp + 31]
"00111111111111100000000000100000",	-- 2688: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 2689: 	addi	%sp, %sp, 33
"01011000000000000000010100000000",	-- 2690: 	jal	sgn.2568
"10101011110111100000000000100001",	-- 2691: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 2692: 	lw	%ra, [%sp + 32]
"10010011110000010000000000011111",	-- 2693: 	lf	%f1, [%sp + 31]
"10110000000111100000000000100000",	-- 2694: 	sf	%f0, [%sp + 32]
"00001100001000000000000000000000",	-- 2695: 	movf	%f0, %f1
"00111111111111100000000000100001",	-- 2696: 	sw	%ra, [%sp + 33]
"10100111110111100000000000100010",	-- 2697: 	addi	%sp, %sp, 34
"01011000000000000000010011101111",	-- 2698: 	jal	fsqr.2530
"10101011110111100000000000100010",	-- 2699: 	subi	%sp, %sp, 34
"00111011110111110000000000100001",	-- 2700: 	lw	%ra, [%sp + 33]
"10010011110000010000000000100000",	-- 2701: 	lf	%f1, [%sp + 32]
"11101100001000000000000000000000",	-- 2702: 	divf	%f0, %f1, %f0
"01010100000000000000101010010010",	-- 2703: 	j	bneq_cont.8971
	-- bneq_else.8970:
"00010100000000000000000000000000",	-- 2704: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2705: 	lhif	%f0, 0.000000
	-- bneq_cont.8971:
"00111011110000010000000000011110",	-- 2706: 	lw	%r1, [%sp + 30]
"00111011110000100000000000000111",	-- 2707: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 2708: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2709: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2710: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 2711: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 2712: 	lf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2713: 	lli	%r1, 2
"00111100001111100000000000100001",	-- 2714: 	sw	%r1, [%sp + 33]
"10110000000111100000000000100010",	-- 2715: 	sf	%f0, [%sp + 34]
"00111111111111100000000000100011",	-- 2716: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 2717: 	addi	%sp, %sp, 36
"01011000000000000000010011100010",	-- 2718: 	jal	fiszero.2526
"10101011110111100000000000100100",	-- 2719: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 2720: 	lw	%ra, [%sp + 35]
"11001100000000100000000000000000",	-- 2721: 	lli	%r2, 0
"00101000001000100000000000010010",	-- 2722: 	bneq	%r1, %r2, bneq_else.8972
"10010011110000000000000000100010",	-- 2723: 	lf	%f0, [%sp + 34]
"00111111111111100000000000100011",	-- 2724: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 2725: 	addi	%sp, %sp, 36
"01011000000000000000010100000000",	-- 2726: 	jal	sgn.2568
"10101011110111100000000000100100",	-- 2727: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 2728: 	lw	%ra, [%sp + 35]
"10010011110000010000000000100010",	-- 2729: 	lf	%f1, [%sp + 34]
"10110000000111100000000000100011",	-- 2730: 	sf	%f0, [%sp + 35]
"00001100001000000000000000000000",	-- 2731: 	movf	%f0, %f1
"00111111111111100000000000100100",	-- 2732: 	sw	%ra, [%sp + 36]
"10100111110111100000000000100101",	-- 2733: 	addi	%sp, %sp, 37
"01011000000000000000010011101111",	-- 2734: 	jal	fsqr.2530
"10101011110111100000000000100101",	-- 2735: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 2736: 	lw	%ra, [%sp + 36]
"10010011110000010000000000100011",	-- 2737: 	lf	%f1, [%sp + 35]
"11101100001000000000000000000000",	-- 2738: 	divf	%f0, %f1, %f0
"01010100000000000000101010110110",	-- 2739: 	j	bneq_cont.8973
	-- bneq_else.8972:
"00010100000000000000000000000000",	-- 2740: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2741: 	lhif	%f0, 0.000000
	-- bneq_cont.8973:
"00111011110000010000000000100001",	-- 2742: 	lw	%r1, [%sp + 33]
"00111011110000100000000000000111",	-- 2743: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 2744: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2745: 	sf	%f0, [%r1 + 0]
"01010100000000000000101011001010",	-- 2746: 	j	bneq_cont.8967
	-- bneq_else.8966:
"11001100000000100000000000000010",	-- 2747: 	lli	%r2, 2
"00101000101000100000000000001110",	-- 2748: 	bneq	%r5, %r2, bneq_else.8974
"11001100000000100000000000000000",	-- 2749: 	lli	%r2, 0
"00111011110001010000000000001110",	-- 2750: 	lw	%r5, [%sp + 14]
"00101000101000100000000000000011",	-- 2751: 	bneq	%r5, %r2, bneq_else.8976
"11001100000000100000000000000001",	-- 2752: 	lli	%r2, 1
"01010100000000000000101011000011",	-- 2753: 	j	bneq_cont.8977
	-- bneq_else.8976:
"11001100000000100000000000000000",	-- 2754: 	lli	%r2, 0
	-- bneq_cont.8977:
"10000100000000110000100000000000",	-- 2755: 	add	%r1, %r0, %r3
"00111111111111100000000000100100",	-- 2756: 	sw	%ra, [%sp + 36]
"10100111110111100000000000100101",	-- 2757: 	addi	%sp, %sp, 37
"01011000000000000000010101001110",	-- 2758: 	jal	vecunit_sgn.2594
"10101011110111100000000000100101",	-- 2759: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 2760: 	lw	%ra, [%sp + 36]
"01010100000000000000101011001010",	-- 2761: 	j	bneq_cont.8975
	-- bneq_else.8974:
	-- bneq_cont.8975:
	-- bneq_cont.8967:
"11001100000000010000000000000000",	-- 2762: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 2763: 	lw	%r2, [%sp + 5]
"00101000010000010000000000000010",	-- 2764: 	bneq	%r2, %r1, bneq_else.8978
"01010100000000000000101011010101",	-- 2765: 	j	bneq_cont.8979
	-- bneq_else.8978:
"00111011110000010000000000000111",	-- 2766: 	lw	%r1, [%sp + 7]
"00111011110000100000000000010110",	-- 2767: 	lw	%r2, [%sp + 22]
"00111111111111100000000000100100",	-- 2768: 	sw	%ra, [%sp + 36]
"10100111110111100000000000100101",	-- 2769: 	addi	%sp, %sp, 37
"01011000000000000000011111110111",	-- 2770: 	jal	rotate_quadratic_matrix.2699
"10101011110111100000000000100101",	-- 2771: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 2772: 	lw	%ra, [%sp + 36]
	-- bneq_cont.8979:
"11001100000000010000000000000001",	-- 2773: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 2774: 	jr	%ra
	-- read_object.2704:
"00111011011000100000000000000010",	-- 2775: 	lw	%r2, [%r27 + 2]
"00111011011000110000000000000001",	-- 2776: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000111100",	-- 2777: 	lli	%r4, 60
"00110000100000010000000000000010",	-- 2778: 	bgt	%r4, %r1, bgt_else.8980
"01001111111000000000000000000000",	-- 2779: 	jr	%ra
	-- bgt_else.8980:
"00111111011111100000000000000000",	-- 2780: 	sw	%r27, [%sp + 0]
"00111100001111100000000000000001",	-- 2781: 	sw	%r1, [%sp + 1]
"00111100011111100000000000000010",	-- 2782: 	sw	%r3, [%sp + 2]
"10000100000000101101100000000000",	-- 2783: 	add	%r27, %r0, %r2
"00111111111111100000000000000011",	-- 2784: 	sw	%ra, [%sp + 3]
"00111011011110100000000000000000",	-- 2785: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000100",	-- 2786: 	addi	%sp, %sp, 4
"01010011010000000000000000000000",	-- 2787: 	jalr	%r26
"10101011110111100000000000000100",	-- 2788: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 2789: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000000",	-- 2790: 	lli	%r2, 0
"00101000001000100000000000000111",	-- 2791: 	bneq	%r1, %r2, bneq_else.8982
"11001100000000010000000000000000",	-- 2792: 	lli	%r1, 0
"00111011110000100000000000000010",	-- 2793: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 2794: 	add	%r1, %r2, %r1
"00111011110000100000000000000001",	-- 2795: 	lw	%r2, [%sp + 1]
"00111100010000010000000000000000",	-- 2796: 	sw	%r2, [%r1 + 0]
"01001111111000000000000000000000",	-- 2797: 	jr	%ra
	-- bneq_else.8982:
"11001100000000010000000000000001",	-- 2798: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 2799: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2800: 	add	%r1, %r2, %r1
"00111011110110110000000000000000",	-- 2801: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 2802: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 2803: 	jr	%r26
	-- read_all_object.2706:
"00111011011110110000000000000001",	-- 2804: 	lw	%r27, [%r27 + 1]
"11001100000000010000000000000000",	-- 2805: 	lli	%r1, 0
"00111011011110100000000000000000",	-- 2806: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 2807: 	jr	%r26
	-- read_net_item.2708:
"00111100001111100000000000000000",	-- 2808: 	sw	%r1, [%sp + 0]
"00111111111111100000000000000001",	-- 2809: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 2810: 	addi	%sp, %sp, 2
"01011000000000000010101000110010",	-- 2811: 	jal	yj_read_int
"10101011110111100000000000000010",	-- 2812: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 2813: 	lw	%ra, [%sp + 1]
"11001100000000101111111111111111",	-- 2814: 	lli	%r2, -1
"11001000000000101111111111111111",	-- 2815: 	lhi	%r2, -1
"00101000001000100000000000000111",	-- 2816: 	bneq	%r1, %r2, bneq_else.8984
"11001100000000010000000000000001",	-- 2817: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 2818: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 2819: 	add	%r1, %r2, %r1
"11001100000000101111111111111111",	-- 2820: 	lli	%r2, -1
"11001000000000101111111111111111",	-- 2821: 	lhi	%r2, -1
"01010100000000000010101000011010",	-- 2822: 	j	yj_create_array
	-- bneq_else.8984:
"11001100000000100000000000000001",	-- 2823: 	lli	%r2, 1
"00111011110000110000000000000000",	-- 2824: 	lw	%r3, [%sp + 0]
"10000100011000100001000000000000",	-- 2825: 	add	%r2, %r3, %r2
"00111100001111100000000000000001",	-- 2826: 	sw	%r1, [%sp + 1]
"10000100000000100000100000000000",	-- 2827: 	add	%r1, %r0, %r2
"00111111111111100000000000000010",	-- 2828: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 2829: 	addi	%sp, %sp, 3
"01011000000000000000101011111000",	-- 2830: 	jal	read_net_item.2708
"10101011110111100000000000000011",	-- 2831: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 2832: 	lw	%ra, [%sp + 2]
"00111011110000100000000000000000",	-- 2833: 	lw	%r2, [%sp + 0]
"10000100001000100001000000000000",	-- 2834: 	add	%r2, %r1, %r2
"00111011110000110000000000000001",	-- 2835: 	lw	%r3, [%sp + 1]
"00111100011000100000000000000000",	-- 2836: 	sw	%r3, [%r2 + 0]
"01001111111000000000000000000000",	-- 2837: 	jr	%ra
	-- read_or_network.2710:
"11001100000000100000000000000000",	-- 2838: 	lli	%r2, 0
"00111100001111100000000000000000",	-- 2839: 	sw	%r1, [%sp + 0]
"10000100000000100000100000000000",	-- 2840: 	add	%r1, %r0, %r2
"00111111111111100000000000000001",	-- 2841: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 2842: 	addi	%sp, %sp, 2
"01011000000000000000101011111000",	-- 2843: 	jal	read_net_item.2708
"10101011110111100000000000000010",	-- 2844: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 2845: 	lw	%ra, [%sp + 1]
"10000100000000010001000000000000",	-- 2846: 	add	%r2, %r0, %r1
"11001100000000010000000000000000",	-- 2847: 	lli	%r1, 0
"10000100010000010000100000000000",	-- 2848: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 2849: 	lw	%r1, [%r1 + 0]
"11001100000000111111111111111111",	-- 2850: 	lli	%r3, -1
"11001000000000111111111111111111",	-- 2851: 	lhi	%r3, -1
"00101000001000110000000000000101",	-- 2852: 	bneq	%r1, %r3, bneq_else.8985
"11001100000000010000000000000001",	-- 2853: 	lli	%r1, 1
"00111011110000110000000000000000",	-- 2854: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 2855: 	add	%r1, %r3, %r1
"01010100000000000010101000011010",	-- 2856: 	j	yj_create_array
	-- bneq_else.8985:
"11001100000000010000000000000001",	-- 2857: 	lli	%r1, 1
"00111011110000110000000000000000",	-- 2858: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 2859: 	add	%r1, %r3, %r1
"00111100010111100000000000000001",	-- 2860: 	sw	%r2, [%sp + 1]
"00111111111111100000000000000010",	-- 2861: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 2862: 	addi	%sp, %sp, 3
"01011000000000000000101100010110",	-- 2863: 	jal	read_or_network.2710
"10101011110111100000000000000011",	-- 2864: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 2865: 	lw	%ra, [%sp + 2]
"00111011110000100000000000000000",	-- 2866: 	lw	%r2, [%sp + 0]
"10000100001000100001000000000000",	-- 2867: 	add	%r2, %r1, %r2
"00111011110000110000000000000001",	-- 2868: 	lw	%r3, [%sp + 1]
"00111100011000100000000000000000",	-- 2869: 	sw	%r3, [%r2 + 0]
"01001111111000000000000000000000",	-- 2870: 	jr	%ra
	-- read_and_network.2712:
"00111011011000100000000000000001",	-- 2871: 	lw	%r2, [%r27 + 1]
"11001100000000110000000000000000",	-- 2872: 	lli	%r3, 0
"00111111011111100000000000000000",	-- 2873: 	sw	%r27, [%sp + 0]
"00111100001111100000000000000001",	-- 2874: 	sw	%r1, [%sp + 1]
"00111100010111100000000000000010",	-- 2875: 	sw	%r2, [%sp + 2]
"10000100000000110000100000000000",	-- 2876: 	add	%r1, %r0, %r3
"00111111111111100000000000000011",	-- 2877: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 2878: 	addi	%sp, %sp, 4
"01011000000000000000101011111000",	-- 2879: 	jal	read_net_item.2708
"10101011110111100000000000000100",	-- 2880: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 2881: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000000",	-- 2882: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 2883: 	add	%r2, %r1, %r2
"00111000010000100000000000000000",	-- 2884: 	lw	%r2, [%r2 + 0]
"11001100000000111111111111111111",	-- 2885: 	lli	%r3, -1
"11001000000000111111111111111111",	-- 2886: 	lhi	%r3, -1
"00101000010000110000000000000010",	-- 2887: 	bneq	%r2, %r3, bneq_else.8986
"01001111111000000000000000000000",	-- 2888: 	jr	%ra
	-- bneq_else.8986:
"00111011110000100000000000000001",	-- 2889: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000010",	-- 2890: 	lw	%r3, [%sp + 2]
"10000100011000100001100000000000",	-- 2891: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 2892: 	sw	%r1, [%r3 + 0]
"11001100000000010000000000000001",	-- 2893: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 2894: 	add	%r1, %r2, %r1
"00111011110110110000000000000000",	-- 2895: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 2896: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 2897: 	jr	%r26
	-- read_parameter.2714:
"00111011011000010000000000000101",	-- 2898: 	lw	%r1, [%r27 + 5]
"00111011011000100000000000000100",	-- 2899: 	lw	%r2, [%r27 + 4]
"00111011011000110000000000000011",	-- 2900: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 2901: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 2902: 	lw	%r5, [%r27 + 1]
"00111100101111100000000000000000",	-- 2903: 	sw	%r5, [%sp + 0]
"00111100011111100000000000000001",	-- 2904: 	sw	%r3, [%sp + 1]
"00111100100111100000000000000010",	-- 2905: 	sw	%r4, [%sp + 2]
"00111100010111100000000000000011",	-- 2906: 	sw	%r2, [%sp + 3]
"10000100000000011101100000000000",	-- 2907: 	add	%r27, %r0, %r1
"00111111111111100000000000000100",	-- 2908: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 2909: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 2910: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 2911: 	jalr	%r26
"10101011110111100000000000000101",	-- 2912: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 2913: 	lw	%ra, [%sp + 4]
"00111011110110110000000000000011",	-- 2914: 	lw	%r27, [%sp + 3]
"00111111111111100000000000000100",	-- 2915: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 2916: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 2917: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 2918: 	jalr	%r26
"10101011110111100000000000000101",	-- 2919: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 2920: 	lw	%ra, [%sp + 4]
"00111011110110110000000000000010",	-- 2921: 	lw	%r27, [%sp + 2]
"00111111111111100000000000000100",	-- 2922: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 2923: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 2924: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 2925: 	jalr	%r26
"10101011110111100000000000000101",	-- 2926: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 2927: 	lw	%ra, [%sp + 4]
"11001100000000010000000000000000",	-- 2928: 	lli	%r1, 0
"00111011110110110000000000000001",	-- 2929: 	lw	%r27, [%sp + 1]
"00111111111111100000000000000100",	-- 2930: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 2931: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 2932: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 2933: 	jalr	%r26
"10101011110111100000000000000101",	-- 2934: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 2935: 	lw	%ra, [%sp + 4]
"11001100000000010000000000000000",	-- 2936: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 2937: 	lli	%r2, 0
"00111100001111100000000000000100",	-- 2938: 	sw	%r1, [%sp + 4]
"10000100000000100000100000000000",	-- 2939: 	add	%r1, %r0, %r2
"00111111111111100000000000000101",	-- 2940: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 2941: 	addi	%sp, %sp, 6
"01011000000000000000101100010110",	-- 2942: 	jal	read_or_network.2710
"10101011110111100000000000000110",	-- 2943: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 2944: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000100",	-- 2945: 	lw	%r2, [%sp + 4]
"00111011110000110000000000000000",	-- 2946: 	lw	%r3, [%sp + 0]
"10000100011000100001000000000000",	-- 2947: 	add	%r2, %r3, %r2
"00111100001000100000000000000000",	-- 2948: 	sw	%r1, [%r2 + 0]
"01001111111000000000000000000000",	-- 2949: 	jr	%ra
	-- solver_rect_surface.2716:
"00111011011001100000000000000001",	-- 2950: 	lw	%r6, [%r27 + 1]
"10000100010000110011100000000000",	-- 2951: 	add	%r7, %r2, %r3
"10010000111000110000000000000000",	-- 2952: 	lf	%f3, [%r7 + 0]
"00111100110111100000000000000000",	-- 2953: 	sw	%r6, [%sp + 0]
"10110000010111100000000000000001",	-- 2954: 	sf	%f2, [%sp + 1]
"00111100101111100000000000000010",	-- 2955: 	sw	%r5, [%sp + 2]
"10110000001111100000000000000011",	-- 2956: 	sf	%f1, [%sp + 3]
"00111100100111100000000000000100",	-- 2957: 	sw	%r4, [%sp + 4]
"10110000000111100000000000000101",	-- 2958: 	sf	%f0, [%sp + 5]
"00111100011111100000000000000110",	-- 2959: 	sw	%r3, [%sp + 6]
"00111100010111100000000000000111",	-- 2960: 	sw	%r2, [%sp + 7]
"00111100001111100000000000001000",	-- 2961: 	sw	%r1, [%sp + 8]
"00001100011000000000000000000000",	-- 2962: 	movf	%f0, %f3
"00111111111111100000000000001001",	-- 2963: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 2964: 	addi	%sp, %sp, 10
"01011000000000000000010011100010",	-- 2965: 	jal	fiszero.2526
"10101011110111100000000000001010",	-- 2966: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 2967: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000000",	-- 2968: 	lli	%r2, 0
"00101000001000100000000001101011",	-- 2969: 	bneq	%r1, %r2, bneq_else.8989
"00111011110000010000000000001000",	-- 2970: 	lw	%r1, [%sp + 8]
"00111111111111100000000000001001",	-- 2971: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 2972: 	addi	%sp, %sp, 10
"01011000000000000000011001100111",	-- 2973: 	jal	o_param_abc.2638
"10101011110111100000000000001010",	-- 2974: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 2975: 	lw	%ra, [%sp + 9]
"00111011110000100000000000001000",	-- 2976: 	lw	%r2, [%sp + 8]
"00111100001111100000000000001001",	-- 2977: 	sw	%r1, [%sp + 9]
"10000100000000100000100000000000",	-- 2978: 	add	%r1, %r0, %r2
"00111111111111100000000000001010",	-- 2979: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 2980: 	addi	%sp, %sp, 11
"01011000000000000000011001010100",	-- 2981: 	jal	o_isinvert.2628
"10101011110111100000000000001011",	-- 2982: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 2983: 	lw	%ra, [%sp + 10]
"00111011110000100000000000000110",	-- 2984: 	lw	%r2, [%sp + 6]
"00111011110000110000000000000111",	-- 2985: 	lw	%r3, [%sp + 7]
"10000100011000100010000000000000",	-- 2986: 	add	%r4, %r3, %r2
"10010000100000000000000000000000",	-- 2987: 	lf	%f0, [%r4 + 0]
"00111100001111100000000000001010",	-- 2988: 	sw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 2989: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 2990: 	addi	%sp, %sp, 12
"01011000000000000000010011011011",	-- 2991: 	jal	fisneg.2524
"10101011110111100000000000001100",	-- 2992: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 2993: 	lw	%ra, [%sp + 11]
"10000100000000010001000000000000",	-- 2994: 	add	%r2, %r0, %r1
"00111011110000010000000000001010",	-- 2995: 	lw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 2996: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 2997: 	addi	%sp, %sp, 12
"01011000000000000000010011110110",	-- 2998: 	jal	xor.2565
"10101011110111100000000000001100",	-- 2999: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3000: 	lw	%ra, [%sp + 11]
"00111011110000100000000000000110",	-- 3001: 	lw	%r2, [%sp + 6]
"00111011110000110000000000001001",	-- 3002: 	lw	%r3, [%sp + 9]
"10000100011000100010000000000000",	-- 3003: 	add	%r4, %r3, %r2
"10010000100000000000000000000000",	-- 3004: 	lf	%f0, [%r4 + 0]
"00111111111111100000000000001011",	-- 3005: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 3006: 	addi	%sp, %sp, 12
"01011000000000000000010100011001",	-- 3007: 	jal	fneg_cond.2570
"10101011110111100000000000001100",	-- 3008: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3009: 	lw	%ra, [%sp + 11]
"10010011110000010000000000000101",	-- 3010: 	lf	%f1, [%sp + 5]
"11100100000000010000000000000000",	-- 3011: 	subf	%f0, %f0, %f1
"00111011110000010000000000000110",	-- 3012: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000111",	-- 3013: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 3014: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3015: 	lf	%f1, [%r1 + 0]
"11101100000000010000000000000000",	-- 3016: 	divf	%f0, %f0, %f1
"00111011110000010000000000000100",	-- 3017: 	lw	%r1, [%sp + 4]
"10000100010000010001100000000000",	-- 3018: 	add	%r3, %r2, %r1
"10010000011000010000000000000000",	-- 3019: 	lf	%f1, [%r3 + 0]
"11101000000000010000100000000000",	-- 3020: 	mulf	%f1, %f0, %f1
"10010011110000100000000000000011",	-- 3021: 	lf	%f2, [%sp + 3]
"11100000001000100000100000000000",	-- 3022: 	addf	%f1, %f1, %f2
"10110000000111100000000000001011",	-- 3023: 	sf	%f0, [%sp + 11]
"00001100001000000000000000000000",	-- 3024: 	movf	%f0, %f1
"00111111111111100000000000001100",	-- 3025: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3026: 	addi	%sp, %sp, 13
"01011000000000000010101001001101",	-- 3027: 	jal	yj_fabs
"10101011110111100000000000001101",	-- 3028: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3029: 	lw	%ra, [%sp + 12]
"00111011110000010000000000000100",	-- 3030: 	lw	%r1, [%sp + 4]
"00111011110000100000000000001001",	-- 3031: 	lw	%r2, [%sp + 9]
"10000100010000010000100000000000",	-- 3032: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3033: 	lf	%f1, [%r1 + 0]
"00111111111111100000000000001100",	-- 3034: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3035: 	addi	%sp, %sp, 13
"01011000000000000000010011110001",	-- 3036: 	jal	fless.2532
"10101011110111100000000000001101",	-- 3037: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3038: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000000",	-- 3039: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3040: 	bneq	%r1, %r2, bneq_else.8990
"11001100000000010000000000000000",	-- 3041: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3042: 	jr	%ra
	-- bneq_else.8990:
"00111011110000010000000000000010",	-- 3043: 	lw	%r1, [%sp + 2]
"00111011110000100000000000000111",	-- 3044: 	lw	%r2, [%sp + 7]
"10000100010000010001000000000000",	-- 3045: 	add	%r2, %r2, %r1
"10010000010000000000000000000000",	-- 3046: 	lf	%f0, [%r2 + 0]
"10010011110000010000000000001011",	-- 3047: 	lf	%f1, [%sp + 11]
"11101000001000000000000000000000",	-- 3048: 	mulf	%f0, %f1, %f0
"10010011110000100000000000000001",	-- 3049: 	lf	%f2, [%sp + 1]
"11100000000000100000000000000000",	-- 3050: 	addf	%f0, %f0, %f2
"00111111111111100000000000001100",	-- 3051: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3052: 	addi	%sp, %sp, 13
"01011000000000000010101001001101",	-- 3053: 	jal	yj_fabs
"10101011110111100000000000001101",	-- 3054: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3055: 	lw	%ra, [%sp + 12]
"00111011110000010000000000000010",	-- 3056: 	lw	%r1, [%sp + 2]
"00111011110000100000000000001001",	-- 3057: 	lw	%r2, [%sp + 9]
"10000100010000010000100000000000",	-- 3058: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3059: 	lf	%f1, [%r1 + 0]
"00111111111111100000000000001100",	-- 3060: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3061: 	addi	%sp, %sp, 13
"01011000000000000000010011110001",	-- 3062: 	jal	fless.2532
"10101011110111100000000000001101",	-- 3063: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3064: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000000",	-- 3065: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3066: 	bneq	%r1, %r2, bneq_else.8991
"11001100000000010000000000000000",	-- 3067: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3068: 	jr	%ra
	-- bneq_else.8991:
"11001100000000010000000000000000",	-- 3069: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 3070: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3071: 	add	%r1, %r2, %r1
"10010011110000000000000000001011",	-- 3072: 	lf	%f0, [%sp + 11]
"10110000000000010000000000000000",	-- 3073: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 3074: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 3075: 	jr	%ra
	-- bneq_else.8989:
"11001100000000010000000000000000",	-- 3076: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3077: 	jr	%ra
	-- solver_rect.2725:
"00111011011110110000000000000001",	-- 3078: 	lw	%r27, [%r27 + 1]
"11001100000000110000000000000000",	-- 3079: 	lli	%r3, 0
"11001100000001000000000000000001",	-- 3080: 	lli	%r4, 1
"11001100000001010000000000000010",	-- 3081: 	lli	%r5, 2
"10110000000111100000000000000000",	-- 3082: 	sf	%f0, [%sp + 0]
"10110000010111100000000000000001",	-- 3083: 	sf	%f2, [%sp + 1]
"10110000001111100000000000000010",	-- 3084: 	sf	%f1, [%sp + 2]
"00111100010111100000000000000011",	-- 3085: 	sw	%r2, [%sp + 3]
"00111100001111100000000000000100",	-- 3086: 	sw	%r1, [%sp + 4]
"00111111011111100000000000000101",	-- 3087: 	sw	%r27, [%sp + 5]
"00111111111111100000000000000110",	-- 3088: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 3089: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 3090: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 3091: 	jalr	%r26
"10101011110111100000000000000111",	-- 3092: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 3093: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 3094: 	lli	%r2, 0
"00101000001000100000000000101001",	-- 3095: 	bneq	%r1, %r2, bneq_else.8992
"11001100000000110000000000000001",	-- 3096: 	lli	%r3, 1
"11001100000001000000000000000010",	-- 3097: 	lli	%r4, 2
"11001100000001010000000000000000",	-- 3098: 	lli	%r5, 0
"10010011110000000000000000000010",	-- 3099: 	lf	%f0, [%sp + 2]
"10010011110000010000000000000001",	-- 3100: 	lf	%f1, [%sp + 1]
"10010011110000100000000000000000",	-- 3101: 	lf	%f2, [%sp + 0]
"00111011110000010000000000000100",	-- 3102: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000011",	-- 3103: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000101",	-- 3104: 	lw	%r27, [%sp + 5]
"00111111111111100000000000000110",	-- 3105: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 3106: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 3107: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 3108: 	jalr	%r26
"10101011110111100000000000000111",	-- 3109: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 3110: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 3111: 	lli	%r2, 0
"00101000001000100000000000010110",	-- 3112: 	bneq	%r1, %r2, bneq_else.8993
"11001100000000110000000000000010",	-- 3113: 	lli	%r3, 2
"11001100000001000000000000000000",	-- 3114: 	lli	%r4, 0
"11001100000001010000000000000001",	-- 3115: 	lli	%r5, 1
"10010011110000000000000000000001",	-- 3116: 	lf	%f0, [%sp + 1]
"10010011110000010000000000000000",	-- 3117: 	lf	%f1, [%sp + 0]
"10010011110000100000000000000010",	-- 3118: 	lf	%f2, [%sp + 2]
"00111011110000010000000000000100",	-- 3119: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000011",	-- 3120: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000101",	-- 3121: 	lw	%r27, [%sp + 5]
"00111111111111100000000000000110",	-- 3122: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 3123: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 3124: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 3125: 	jalr	%r26
"10101011110111100000000000000111",	-- 3126: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 3127: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 3128: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3129: 	bneq	%r1, %r2, bneq_else.8994
"11001100000000010000000000000000",	-- 3130: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3131: 	jr	%ra
	-- bneq_else.8994:
"11001100000000010000000000000011",	-- 3132: 	lli	%r1, 3
"01001111111000000000000000000000",	-- 3133: 	jr	%ra
	-- bneq_else.8993:
"11001100000000010000000000000010",	-- 3134: 	lli	%r1, 2
"01001111111000000000000000000000",	-- 3135: 	jr	%ra
	-- bneq_else.8992:
"11001100000000010000000000000001",	-- 3136: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 3137: 	jr	%ra
	-- solver_surface.2731:
"00111011011000110000000000000001",	-- 3138: 	lw	%r3, [%r27 + 1]
"00111100011111100000000000000000",	-- 3139: 	sw	%r3, [%sp + 0]
"10110000010111100000000000000001",	-- 3140: 	sf	%f2, [%sp + 1]
"10110000001111100000000000000010",	-- 3141: 	sf	%f1, [%sp + 2]
"10110000000111100000000000000011",	-- 3142: 	sf	%f0, [%sp + 3]
"00111100010111100000000000000100",	-- 3143: 	sw	%r2, [%sp + 4]
"00111111111111100000000000000101",	-- 3144: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 3145: 	addi	%sp, %sp, 6
"01011000000000000000011001100111",	-- 3146: 	jal	o_param_abc.2638
"10101011110111100000000000000110",	-- 3147: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 3148: 	lw	%ra, [%sp + 5]
"10000100000000010001000000000000",	-- 3149: 	add	%r2, %r0, %r1
"00111011110000010000000000000100",	-- 3150: 	lw	%r1, [%sp + 4]
"00111100010111100000000000000101",	-- 3151: 	sw	%r2, [%sp + 5]
"00111111111111100000000000000110",	-- 3152: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 3153: 	addi	%sp, %sp, 7
"01011000000000000000010110100101",	-- 3154: 	jal	veciprod.2597
"10101011110111100000000000000111",	-- 3155: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 3156: 	lw	%ra, [%sp + 6]
"10110000000111100000000000000110",	-- 3157: 	sf	%f0, [%sp + 6]
"00111111111111100000000000000111",	-- 3158: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 3159: 	addi	%sp, %sp, 8
"01011000000000000000010011010100",	-- 3160: 	jal	fispos.2522
"10101011110111100000000000001000",	-- 3161: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 3162: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000000",	-- 3163: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3164: 	bneq	%r1, %r2, bneq_else.8995
"11001100000000010000000000000000",	-- 3165: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3166: 	jr	%ra
	-- bneq_else.8995:
"11001100000000010000000000000000",	-- 3167: 	lli	%r1, 0
"10010011110000000000000000000011",	-- 3168: 	lf	%f0, [%sp + 3]
"10010011110000010000000000000010",	-- 3169: 	lf	%f1, [%sp + 2]
"10010011110000100000000000000001",	-- 3170: 	lf	%f2, [%sp + 1]
"00111011110000100000000000000101",	-- 3171: 	lw	%r2, [%sp + 5]
"00111100001111100000000000000111",	-- 3172: 	sw	%r1, [%sp + 7]
"10000100000000100000100000000000",	-- 3173: 	add	%r1, %r0, %r2
"00111111111111100000000000001000",	-- 3174: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 3175: 	addi	%sp, %sp, 9
"01011000000000000000010110111101",	-- 3176: 	jal	veciprod2.2600
"10101011110111100000000000001001",	-- 3177: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 3178: 	lw	%ra, [%sp + 8]
"00111111111111100000000000001000",	-- 3179: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 3180: 	addi	%sp, %sp, 9
"01011000000000000010101001001111",	-- 3181: 	jal	yj_fneg
"10101011110111100000000000001001",	-- 3182: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 3183: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000110",	-- 3184: 	lf	%f1, [%sp + 6]
"11101100000000010000000000000000",	-- 3185: 	divf	%f0, %f0, %f1
"00111011110000010000000000000111",	-- 3186: 	lw	%r1, [%sp + 7]
"00111011110000100000000000000000",	-- 3187: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3188: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 3189: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 3190: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 3191: 	jr	%ra
	-- quadratic.2737:
"10110000000111100000000000000000",	-- 3192: 	sf	%f0, [%sp + 0]
"10110000010111100000000000000001",	-- 3193: 	sf	%f2, [%sp + 1]
"10110000001111100000000000000010",	-- 3194: 	sf	%f1, [%sp + 2]
"00111100001111100000000000000011",	-- 3195: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 3196: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 3197: 	addi	%sp, %sp, 5
"01011000000000000000010011101111",	-- 3198: 	jal	fsqr.2530
"10101011110111100000000000000101",	-- 3199: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 3200: 	lw	%ra, [%sp + 4]
"00111011110000010000000000000011",	-- 3201: 	lw	%r1, [%sp + 3]
"10110000000111100000000000000100",	-- 3202: 	sf	%f0, [%sp + 4]
"00111111111111100000000000000101",	-- 3203: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 3204: 	addi	%sp, %sp, 6
"01011000000000000000011001011000",	-- 3205: 	jal	o_param_a.2632
"10101011110111100000000000000110",	-- 3206: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 3207: 	lw	%ra, [%sp + 5]
"10010011110000010000000000000100",	-- 3208: 	lf	%f1, [%sp + 4]
"11101000001000000000000000000000",	-- 3209: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000010",	-- 3210: 	lf	%f1, [%sp + 2]
"10110000000111100000000000000101",	-- 3211: 	sf	%f0, [%sp + 5]
"00001100001000000000000000000000",	-- 3212: 	movf	%f0, %f1
"00111111111111100000000000000110",	-- 3213: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 3214: 	addi	%sp, %sp, 7
"01011000000000000000010011101111",	-- 3215: 	jal	fsqr.2530
"10101011110111100000000000000111",	-- 3216: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 3217: 	lw	%ra, [%sp + 6]
"00111011110000010000000000000011",	-- 3218: 	lw	%r1, [%sp + 3]
"10110000000111100000000000000110",	-- 3219: 	sf	%f0, [%sp + 6]
"00111111111111100000000000000111",	-- 3220: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 3221: 	addi	%sp, %sp, 8
"01011000000000000000011001011101",	-- 3222: 	jal	o_param_b.2634
"10101011110111100000000000001000",	-- 3223: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 3224: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000110",	-- 3225: 	lf	%f1, [%sp + 6]
"11101000001000000000000000000000",	-- 3226: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000101",	-- 3227: 	lf	%f1, [%sp + 5]
"11100000001000000000000000000000",	-- 3228: 	addf	%f0, %f1, %f0
"10010011110000010000000000000001",	-- 3229: 	lf	%f1, [%sp + 1]
"10110000000111100000000000000111",	-- 3230: 	sf	%f0, [%sp + 7]
"00001100001000000000000000000000",	-- 3231: 	movf	%f0, %f1
"00111111111111100000000000001000",	-- 3232: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 3233: 	addi	%sp, %sp, 9
"01011000000000000000010011101111",	-- 3234: 	jal	fsqr.2530
"10101011110111100000000000001001",	-- 3235: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 3236: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000011",	-- 3237: 	lw	%r1, [%sp + 3]
"10110000000111100000000000001000",	-- 3238: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 3239: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 3240: 	addi	%sp, %sp, 10
"01011000000000000000011001100010",	-- 3241: 	jal	o_param_c.2636
"10101011110111100000000000001010",	-- 3242: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 3243: 	lw	%ra, [%sp + 9]
"10010011110000010000000000001000",	-- 3244: 	lf	%f1, [%sp + 8]
"11101000001000000000000000000000",	-- 3245: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000111",	-- 3246: 	lf	%f1, [%sp + 7]
"11100000001000000000000000000000",	-- 3247: 	addf	%f0, %f1, %f0
"00111011110000010000000000000011",	-- 3248: 	lw	%r1, [%sp + 3]
"10110000000111100000000000001001",	-- 3249: 	sf	%f0, [%sp + 9]
"00111111111111100000000000001010",	-- 3250: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 3251: 	addi	%sp, %sp, 11
"01011000000000000000011001010110",	-- 3252: 	jal	o_isrot.2630
"10101011110111100000000000001011",	-- 3253: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 3254: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 3255: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3256: 	bneq	%r1, %r2, bneq_else.8996
"10010011110000000000000000001001",	-- 3257: 	lf	%f0, [%sp + 9]
"01001111111000000000000000000000",	-- 3258: 	jr	%ra
	-- bneq_else.8996:
"10010011110000000000000000000001",	-- 3259: 	lf	%f0, [%sp + 1]
"10010011110000010000000000000010",	-- 3260: 	lf	%f1, [%sp + 2]
"11101000001000000001000000000000",	-- 3261: 	mulf	%f2, %f1, %f0
"00111011110000010000000000000011",	-- 3262: 	lw	%r1, [%sp + 3]
"10110000010111100000000000001010",	-- 3263: 	sf	%f2, [%sp + 10]
"00111111111111100000000000001011",	-- 3264: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 3265: 	addi	%sp, %sp, 12
"01011000000000000000011010010001",	-- 3266: 	jal	o_param_r1.2656
"10101011110111100000000000001100",	-- 3267: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3268: 	lw	%ra, [%sp + 11]
"10010011110000010000000000001010",	-- 3269: 	lf	%f1, [%sp + 10]
"11101000001000000000000000000000",	-- 3270: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001001",	-- 3271: 	lf	%f1, [%sp + 9]
"11100000001000000000000000000000",	-- 3272: 	addf	%f0, %f1, %f0
"10010011110000010000000000000000",	-- 3273: 	lf	%f1, [%sp + 0]
"10010011110000100000000000000001",	-- 3274: 	lf	%f2, [%sp + 1]
"11101000010000010001000000000000",	-- 3275: 	mulf	%f2, %f2, %f1
"00111011110000010000000000000011",	-- 3276: 	lw	%r1, [%sp + 3]
"10110000000111100000000000001011",	-- 3277: 	sf	%f0, [%sp + 11]
"10110000010111100000000000001100",	-- 3278: 	sf	%f2, [%sp + 12]
"00111111111111100000000000001101",	-- 3279: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 3280: 	addi	%sp, %sp, 14
"01011000000000000000011010010110",	-- 3281: 	jal	o_param_r2.2658
"10101011110111100000000000001110",	-- 3282: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 3283: 	lw	%ra, [%sp + 13]
"10010011110000010000000000001100",	-- 3284: 	lf	%f1, [%sp + 12]
"11101000001000000000000000000000",	-- 3285: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001011",	-- 3286: 	lf	%f1, [%sp + 11]
"11100000001000000000000000000000",	-- 3287: 	addf	%f0, %f1, %f0
"10010011110000010000000000000010",	-- 3288: 	lf	%f1, [%sp + 2]
"10010011110000100000000000000000",	-- 3289: 	lf	%f2, [%sp + 0]
"11101000010000010000100000000000",	-- 3290: 	mulf	%f1, %f2, %f1
"00111011110000010000000000000011",	-- 3291: 	lw	%r1, [%sp + 3]
"10110000000111100000000000001101",	-- 3292: 	sf	%f0, [%sp + 13]
"10110000001111100000000000001110",	-- 3293: 	sf	%f1, [%sp + 14]
"00111111111111100000000000001111",	-- 3294: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 3295: 	addi	%sp, %sp, 16
"01011000000000000000011010011011",	-- 3296: 	jal	o_param_r3.2660
"10101011110111100000000000010000",	-- 3297: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 3298: 	lw	%ra, [%sp + 15]
"10010011110000010000000000001110",	-- 3299: 	lf	%f1, [%sp + 14]
"11101000001000000000000000000000",	-- 3300: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001101",	-- 3301: 	lf	%f1, [%sp + 13]
"11100000001000000000000000000000",	-- 3302: 	addf	%f0, %f1, %f0
"01001111111000000000000000000000",	-- 3303: 	jr	%ra
	-- bilinear.2742:
"11101000000000110011000000000000",	-- 3304: 	mulf	%f6, %f0, %f3
"10110000011111100000000000000000",	-- 3305: 	sf	%f3, [%sp + 0]
"10110000000111100000000000000001",	-- 3306: 	sf	%f0, [%sp + 1]
"10110000101111100000000000000010",	-- 3307: 	sf	%f5, [%sp + 2]
"10110000010111100000000000000011",	-- 3308: 	sf	%f2, [%sp + 3]
"00111100001111100000000000000100",	-- 3309: 	sw	%r1, [%sp + 4]
"10110000100111100000000000000101",	-- 3310: 	sf	%f4, [%sp + 5]
"10110000001111100000000000000110",	-- 3311: 	sf	%f1, [%sp + 6]
"10110000110111100000000000000111",	-- 3312: 	sf	%f6, [%sp + 7]
"00111111111111100000000000001000",	-- 3313: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 3314: 	addi	%sp, %sp, 9
"01011000000000000000011001011000",	-- 3315: 	jal	o_param_a.2632
"10101011110111100000000000001001",	-- 3316: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 3317: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000111",	-- 3318: 	lf	%f1, [%sp + 7]
"11101000001000000000000000000000",	-- 3319: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000101",	-- 3320: 	lf	%f1, [%sp + 5]
"10010011110000100000000000000110",	-- 3321: 	lf	%f2, [%sp + 6]
"11101000010000010001100000000000",	-- 3322: 	mulf	%f3, %f2, %f1
"00111011110000010000000000000100",	-- 3323: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001000",	-- 3324: 	sf	%f0, [%sp + 8]
"10110000011111100000000000001001",	-- 3325: 	sf	%f3, [%sp + 9]
"00111111111111100000000000001010",	-- 3326: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 3327: 	addi	%sp, %sp, 11
"01011000000000000000011001011101",	-- 3328: 	jal	o_param_b.2634
"10101011110111100000000000001011",	-- 3329: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 3330: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 3331: 	lf	%f1, [%sp + 9]
"11101000001000000000000000000000",	-- 3332: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001000",	-- 3333: 	lf	%f1, [%sp + 8]
"11100000001000000000000000000000",	-- 3334: 	addf	%f0, %f1, %f0
"10010011110000010000000000000010",	-- 3335: 	lf	%f1, [%sp + 2]
"10010011110000100000000000000011",	-- 3336: 	lf	%f2, [%sp + 3]
"11101000010000010001100000000000",	-- 3337: 	mulf	%f3, %f2, %f1
"00111011110000010000000000000100",	-- 3338: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001010",	-- 3339: 	sf	%f0, [%sp + 10]
"10110000011111100000000000001011",	-- 3340: 	sf	%f3, [%sp + 11]
"00111111111111100000000000001100",	-- 3341: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3342: 	addi	%sp, %sp, 13
"01011000000000000000011001100010",	-- 3343: 	jal	o_param_c.2636
"10101011110111100000000000001101",	-- 3344: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3345: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001011",	-- 3346: 	lf	%f1, [%sp + 11]
"11101000001000000000000000000000",	-- 3347: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001010",	-- 3348: 	lf	%f1, [%sp + 10]
"11100000001000000000000000000000",	-- 3349: 	addf	%f0, %f1, %f0
"00111011110000010000000000000100",	-- 3350: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001100",	-- 3351: 	sf	%f0, [%sp + 12]
"00111111111111100000000000001101",	-- 3352: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 3353: 	addi	%sp, %sp, 14
"01011000000000000000011001010110",	-- 3354: 	jal	o_isrot.2630
"10101011110111100000000000001110",	-- 3355: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 3356: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 3357: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3358: 	bneq	%r1, %r2, bneq_else.8997
"10010011110000000000000000001100",	-- 3359: 	lf	%f0, [%sp + 12]
"01001111111000000000000000000000",	-- 3360: 	jr	%ra
	-- bneq_else.8997:
"10010011110000000000000000000101",	-- 3361: 	lf	%f0, [%sp + 5]
"10010011110000010000000000000011",	-- 3362: 	lf	%f1, [%sp + 3]
"11101000001000000001000000000000",	-- 3363: 	mulf	%f2, %f1, %f0
"10010011110000110000000000000010",	-- 3364: 	lf	%f3, [%sp + 2]
"10010011110001000000000000000110",	-- 3365: 	lf	%f4, [%sp + 6]
"11101000100000110010100000000000",	-- 3366: 	mulf	%f5, %f4, %f3
"11100000010001010001000000000000",	-- 3367: 	addf	%f2, %f2, %f5
"00111011110000010000000000000100",	-- 3368: 	lw	%r1, [%sp + 4]
"10110000010111100000000000001101",	-- 3369: 	sf	%f2, [%sp + 13]
"00111111111111100000000000001110",	-- 3370: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 3371: 	addi	%sp, %sp, 15
"01011000000000000000011010010001",	-- 3372: 	jal	o_param_r1.2656
"10101011110111100000000000001111",	-- 3373: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 3374: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001101",	-- 3375: 	lf	%f1, [%sp + 13]
"11101000001000000000000000000000",	-- 3376: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000010",	-- 3377: 	lf	%f1, [%sp + 2]
"10010011110000100000000000000001",	-- 3378: 	lf	%f2, [%sp + 1]
"11101000010000010000100000000000",	-- 3379: 	mulf	%f1, %f2, %f1
"10010011110000110000000000000000",	-- 3380: 	lf	%f3, [%sp + 0]
"10010011110001000000000000000011",	-- 3381: 	lf	%f4, [%sp + 3]
"11101000100000110010000000000000",	-- 3382: 	mulf	%f4, %f4, %f3
"11100000001001000000100000000000",	-- 3383: 	addf	%f1, %f1, %f4
"00111011110000010000000000000100",	-- 3384: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001110",	-- 3385: 	sf	%f0, [%sp + 14]
"10110000001111100000000000001111",	-- 3386: 	sf	%f1, [%sp + 15]
"00111111111111100000000000010000",	-- 3387: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 3388: 	addi	%sp, %sp, 17
"01011000000000000000011010010110",	-- 3389: 	jal	o_param_r2.2658
"10101011110111100000000000010001",	-- 3390: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 3391: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001111",	-- 3392: 	lf	%f1, [%sp + 15]
"11101000001000000000000000000000",	-- 3393: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001110",	-- 3394: 	lf	%f1, [%sp + 14]
"11100000001000000000000000000000",	-- 3395: 	addf	%f0, %f1, %f0
"10010011110000010000000000000101",	-- 3396: 	lf	%f1, [%sp + 5]
"10010011110000100000000000000001",	-- 3397: 	lf	%f2, [%sp + 1]
"11101000010000010000100000000000",	-- 3398: 	mulf	%f1, %f2, %f1
"10010011110000100000000000000000",	-- 3399: 	lf	%f2, [%sp + 0]
"10010011110000110000000000000110",	-- 3400: 	lf	%f3, [%sp + 6]
"11101000011000100001000000000000",	-- 3401: 	mulf	%f2, %f3, %f2
"11100000001000100000100000000000",	-- 3402: 	addf	%f1, %f1, %f2
"00111011110000010000000000000100",	-- 3403: 	lw	%r1, [%sp + 4]
"10110000000111100000000000010000",	-- 3404: 	sf	%f0, [%sp + 16]
"10110000001111100000000000010001",	-- 3405: 	sf	%f1, [%sp + 17]
"00111111111111100000000000010010",	-- 3406: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 3407: 	addi	%sp, %sp, 19
"01011000000000000000011010011011",	-- 3408: 	jal	o_param_r3.2660
"10101011110111100000000000010011",	-- 3409: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 3410: 	lw	%ra, [%sp + 18]
"10010011110000010000000000010001",	-- 3411: 	lf	%f1, [%sp + 17]
"11101000001000000000000000000000",	-- 3412: 	mulf	%f0, %f1, %f0
"10010011110000010000000000010000",	-- 3413: 	lf	%f1, [%sp + 16]
"11100000001000000000000000000000",	-- 3414: 	addf	%f0, %f1, %f0
"00111111111111100000000000010010",	-- 3415: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 3416: 	addi	%sp, %sp, 19
"01011000000000000000010011101011",	-- 3417: 	jal	fhalf.2528
"10101011110111100000000000010011",	-- 3418: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 3419: 	lw	%ra, [%sp + 18]
"10010011110000010000000000001100",	-- 3420: 	lf	%f1, [%sp + 12]
"11100000001000000000000000000000",	-- 3421: 	addf	%f0, %f1, %f0
"01001111111000000000000000000000",	-- 3422: 	jr	%ra
	-- solver_second.2750:
"00111011011000110000000000000001",	-- 3423: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 3424: 	lli	%r4, 0
"10000100010001000010000000000000",	-- 3425: 	add	%r4, %r2, %r4
"10010000100000110000000000000000",	-- 3426: 	lf	%f3, [%r4 + 0]
"11001100000001000000000000000001",	-- 3427: 	lli	%r4, 1
"10000100010001000010000000000000",	-- 3428: 	add	%r4, %r2, %r4
"10010000100001000000000000000000",	-- 3429: 	lf	%f4, [%r4 + 0]
"11001100000001000000000000000010",	-- 3430: 	lli	%r4, 2
"10000100010001000010000000000000",	-- 3431: 	add	%r4, %r2, %r4
"10010000100001010000000000000000",	-- 3432: 	lf	%f5, [%r4 + 0]
"00111100011111100000000000000000",	-- 3433: 	sw	%r3, [%sp + 0]
"10110000010111100000000000000001",	-- 3434: 	sf	%f2, [%sp + 1]
"10110000001111100000000000000010",	-- 3435: 	sf	%f1, [%sp + 2]
"10110000000111100000000000000011",	-- 3436: 	sf	%f0, [%sp + 3]
"00111100001111100000000000000100",	-- 3437: 	sw	%r1, [%sp + 4]
"00111100010111100000000000000101",	-- 3438: 	sw	%r2, [%sp + 5]
"00001100101000100000000000000000",	-- 3439: 	movf	%f2, %f5
"00001100100000010000000000000000",	-- 3440: 	movf	%f1, %f4
"00001100011000000000000000000000",	-- 3441: 	movf	%f0, %f3
"00111111111111100000000000000110",	-- 3442: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 3443: 	addi	%sp, %sp, 7
"01011000000000000000110001111000",	-- 3444: 	jal	quadratic.2737
"10101011110111100000000000000111",	-- 3445: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 3446: 	lw	%ra, [%sp + 6]
"10110000000111100000000000000110",	-- 3447: 	sf	%f0, [%sp + 6]
"00111111111111100000000000000111",	-- 3448: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 3449: 	addi	%sp, %sp, 8
"01011000000000000000010011100010",	-- 3450: 	jal	fiszero.2526
"10101011110111100000000000001000",	-- 3451: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 3452: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000000",	-- 3453: 	lli	%r2, 0
"00101000001000100000000001100111",	-- 3454: 	bneq	%r1, %r2, bneq_else.8998
"11001100000000010000000000000000",	-- 3455: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 3456: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 3457: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3458: 	lf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 3459: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 3460: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3461: 	lf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 3462: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 3463: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 3464: 	lf	%f2, [%r1 + 0]
"10010011110000110000000000000011",	-- 3465: 	lf	%f3, [%sp + 3]
"10010011110001000000000000000010",	-- 3466: 	lf	%f4, [%sp + 2]
"10010011110001010000000000000001",	-- 3467: 	lf	%f5, [%sp + 1]
"00111011110000010000000000000100",	-- 3468: 	lw	%r1, [%sp + 4]
"00111111111111100000000000000111",	-- 3469: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 3470: 	addi	%sp, %sp, 8
"01011000000000000000110011101000",	-- 3471: 	jal	bilinear.2742
"10101011110111100000000000001000",	-- 3472: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 3473: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000011",	-- 3474: 	lf	%f1, [%sp + 3]
"10010011110000100000000000000010",	-- 3475: 	lf	%f2, [%sp + 2]
"10010011110000110000000000000001",	-- 3476: 	lf	%f3, [%sp + 1]
"00111011110000010000000000000100",	-- 3477: 	lw	%r1, [%sp + 4]
"10110000000111100000000000000111",	-- 3478: 	sf	%f0, [%sp + 7]
"00001100001000000000000000000000",	-- 3479: 	movf	%f0, %f1
"00001100010000010000000000000000",	-- 3480: 	movf	%f1, %f2
"00001100011000100000000000000000",	-- 3481: 	movf	%f2, %f3
"00111111111111100000000000001000",	-- 3482: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 3483: 	addi	%sp, %sp, 9
"01011000000000000000110001111000",	-- 3484: 	jal	quadratic.2737
"10101011110111100000000000001001",	-- 3485: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 3486: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000100",	-- 3487: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001000",	-- 3488: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 3489: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 3490: 	addi	%sp, %sp, 10
"01011000000000000000011001010000",	-- 3491: 	jal	o_form.2624
"10101011110111100000000000001010",	-- 3492: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 3493: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000011",	-- 3494: 	lli	%r2, 3
"00101000001000100000000000000110",	-- 3495: 	bneq	%r1, %r2, bneq_else.8999
"00010100000000000000000000000000",	-- 3496: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 3497: 	lhif	%f0, 1.000000
"10010011110000010000000000001000",	-- 3498: 	lf	%f1, [%sp + 8]
"11100100001000000000000000000000",	-- 3499: 	subf	%f0, %f1, %f0
"01010100000000000000110110101110",	-- 3500: 	j	bneq_cont.9000
	-- bneq_else.8999:
"10010011110000000000000000001000",	-- 3501: 	lf	%f0, [%sp + 8]
	-- bneq_cont.9000:
"10010011110000010000000000000111",	-- 3502: 	lf	%f1, [%sp + 7]
"10110000000111100000000000001001",	-- 3503: 	sf	%f0, [%sp + 9]
"00001100001000000000000000000000",	-- 3504: 	movf	%f0, %f1
"00111111111111100000000000001010",	-- 3505: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 3506: 	addi	%sp, %sp, 11
"01011000000000000000010011101111",	-- 3507: 	jal	fsqr.2530
"10101011110111100000000000001011",	-- 3508: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 3509: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 3510: 	lf	%f1, [%sp + 9]
"10010011110000100000000000000110",	-- 3511: 	lf	%f2, [%sp + 6]
"11101000010000010000100000000000",	-- 3512: 	mulf	%f1, %f2, %f1
"11100100000000010000000000000000",	-- 3513: 	subf	%f0, %f0, %f1
"10110000000111100000000000001010",	-- 3514: 	sf	%f0, [%sp + 10]
"00111111111111100000000000001011",	-- 3515: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 3516: 	addi	%sp, %sp, 12
"01011000000000000000010011010100",	-- 3517: 	jal	fispos.2522
"10101011110111100000000000001100",	-- 3518: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3519: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 3520: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3521: 	bneq	%r1, %r2, bneq_else.9001
"11001100000000010000000000000000",	-- 3522: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3523: 	jr	%ra
	-- bneq_else.9001:
"10010011110000000000000000001010",	-- 3524: 	lf	%f0, [%sp + 10]
"00111111111111100000000000001011",	-- 3525: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 3526: 	addi	%sp, %sp, 12
"01011000000000000010101000101110",	-- 3527: 	jal	yj_sqrt
"10101011110111100000000000001100",	-- 3528: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3529: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000100",	-- 3530: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001011",	-- 3531: 	sf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 3532: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3533: 	addi	%sp, %sp, 13
"01011000000000000000011001010100",	-- 3534: 	jal	o_isinvert.2628
"10101011110111100000000000001101",	-- 3535: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3536: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000000",	-- 3537: 	lli	%r2, 0
"00101000001000100000000000001000",	-- 3538: 	bneq	%r1, %r2, bneq_else.9002
"10010011110000000000000000001011",	-- 3539: 	lf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 3540: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3541: 	addi	%sp, %sp, 13
"01011000000000000010101001001111",	-- 3542: 	jal	yj_fneg
"10101011110111100000000000001101",	-- 3543: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3544: 	lw	%ra, [%sp + 12]
"01010100000000000000110111011011",	-- 3545: 	j	bneq_cont.9003
	-- bneq_else.9002:
"10010011110000000000000000001011",	-- 3546: 	lf	%f0, [%sp + 11]
	-- bneq_cont.9003:
"11001100000000010000000000000000",	-- 3547: 	lli	%r1, 0
"10010011110000010000000000000111",	-- 3548: 	lf	%f1, [%sp + 7]
"11100100000000010000000000000000",	-- 3549: 	subf	%f0, %f0, %f1
"10010011110000010000000000000110",	-- 3550: 	lf	%f1, [%sp + 6]
"11101100000000010000000000000000",	-- 3551: 	divf	%f0, %f0, %f1
"00111011110000100000000000000000",	-- 3552: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3553: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 3554: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 3555: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 3556: 	jr	%ra
	-- bneq_else.8998:
"11001100000000010000000000000000",	-- 3557: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3558: 	jr	%ra
	-- solver.2756:
"00111011011001000000000000000100",	-- 3559: 	lw	%r4, [%r27 + 4]
"00111011011001010000000000000011",	-- 3560: 	lw	%r5, [%r27 + 3]
"00111011011001100000000000000010",	-- 3561: 	lw	%r6, [%r27 + 2]
"00111011011001110000000000000001",	-- 3562: 	lw	%r7, [%r27 + 1]
"10000100111000010000100000000000",	-- 3563: 	add	%r1, %r7, %r1
"00111000001000010000000000000000",	-- 3564: 	lw	%r1, [%r1 + 0]
"11001100000001110000000000000000",	-- 3565: 	lli	%r7, 0
"10000100011001110011100000000000",	-- 3566: 	add	%r7, %r3, %r7
"10010000111000000000000000000000",	-- 3567: 	lf	%f0, [%r7 + 0]
"00111100101111100000000000000000",	-- 3568: 	sw	%r5, [%sp + 0]
"00111100100111100000000000000001",	-- 3569: 	sw	%r4, [%sp + 1]
"00111100010111100000000000000010",	-- 3570: 	sw	%r2, [%sp + 2]
"00111100110111100000000000000011",	-- 3571: 	sw	%r6, [%sp + 3]
"00111100001111100000000000000100",	-- 3572: 	sw	%r1, [%sp + 4]
"00111100011111100000000000000101",	-- 3573: 	sw	%r3, [%sp + 5]
"10110000000111100000000000000110",	-- 3574: 	sf	%f0, [%sp + 6]
"00111111111111100000000000000111",	-- 3575: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 3576: 	addi	%sp, %sp, 8
"01011000000000000000011001101001",	-- 3577: 	jal	o_param_x.2640
"10101011110111100000000000001000",	-- 3578: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 3579: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000110",	-- 3580: 	lf	%f1, [%sp + 6]
"11100100001000000000000000000000",	-- 3581: 	subf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 3582: 	lli	%r1, 1
"00111011110000100000000000000101",	-- 3583: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 3584: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3585: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000100",	-- 3586: 	lw	%r1, [%sp + 4]
"10110000000111100000000000000111",	-- 3587: 	sf	%f0, [%sp + 7]
"10110000001111100000000000001000",	-- 3588: 	sf	%f1, [%sp + 8]
"00111111111111100000000000001001",	-- 3589: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 3590: 	addi	%sp, %sp, 10
"01011000000000000000011001101110",	-- 3591: 	jal	o_param_y.2642
"10101011110111100000000000001010",	-- 3592: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 3593: 	lw	%ra, [%sp + 9]
"10010011110000010000000000001000",	-- 3594: 	lf	%f1, [%sp + 8]
"11100100001000000000000000000000",	-- 3595: 	subf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 3596: 	lli	%r1, 2
"00111011110000100000000000000101",	-- 3597: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 3598: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3599: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000100",	-- 3600: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001001",	-- 3601: 	sf	%f0, [%sp + 9]
"10110000001111100000000000001010",	-- 3602: 	sf	%f1, [%sp + 10]
"00111111111111100000000000001011",	-- 3603: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 3604: 	addi	%sp, %sp, 12
"01011000000000000000011001110011",	-- 3605: 	jal	o_param_z.2644
"10101011110111100000000000001100",	-- 3606: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3607: 	lw	%ra, [%sp + 11]
"10010011110000010000000000001010",	-- 3608: 	lf	%f1, [%sp + 10]
"11100100001000000000000000000000",	-- 3609: 	subf	%f0, %f1, %f0
"00111011110000010000000000000100",	-- 3610: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001011",	-- 3611: 	sf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 3612: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3613: 	addi	%sp, %sp, 13
"01011000000000000000011001010000",	-- 3614: 	jal	o_form.2624
"10101011110111100000000000001101",	-- 3615: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3616: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000001",	-- 3617: 	lli	%r2, 1
"00101000001000100000000000001001",	-- 3618: 	bneq	%r1, %r2, bneq_else.9004
"10010011110000000000000000000111",	-- 3619: 	lf	%f0, [%sp + 7]
"10010011110000010000000000001001",	-- 3620: 	lf	%f1, [%sp + 9]
"10010011110000100000000000001011",	-- 3621: 	lf	%f2, [%sp + 11]
"00111011110000010000000000000100",	-- 3622: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000010",	-- 3623: 	lw	%r2, [%sp + 2]
"00111011110110110000000000000011",	-- 3624: 	lw	%r27, [%sp + 3]
"00111011011110100000000000000000",	-- 3625: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 3626: 	jr	%r26
	-- bneq_else.9004:
"11001100000000100000000000000010",	-- 3627: 	lli	%r2, 2
"00101000001000100000000000001001",	-- 3628: 	bneq	%r1, %r2, bneq_else.9005
"10010011110000000000000000000111",	-- 3629: 	lf	%f0, [%sp + 7]
"10010011110000010000000000001001",	-- 3630: 	lf	%f1, [%sp + 9]
"10010011110000100000000000001011",	-- 3631: 	lf	%f2, [%sp + 11]
"00111011110000010000000000000100",	-- 3632: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000010",	-- 3633: 	lw	%r2, [%sp + 2]
"00111011110110110000000000000001",	-- 3634: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 3635: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 3636: 	jr	%r26
	-- bneq_else.9005:
"10010011110000000000000000000111",	-- 3637: 	lf	%f0, [%sp + 7]
"10010011110000010000000000001001",	-- 3638: 	lf	%f1, [%sp + 9]
"10010011110000100000000000001011",	-- 3639: 	lf	%f2, [%sp + 11]
"00111011110000010000000000000100",	-- 3640: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000010",	-- 3641: 	lw	%r2, [%sp + 2]
"00111011110110110000000000000000",	-- 3642: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 3643: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 3644: 	jr	%r26
	-- solver_rect_fast.2760:
"00111011011001000000000000000001",	-- 3645: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 3646: 	lli	%r5, 0
"10000100011001010010100000000000",	-- 3647: 	add	%r5, %r3, %r5
"10010000101000110000000000000000",	-- 3648: 	lf	%f3, [%r5 + 0]
"11100100011000000001100000000000",	-- 3649: 	subf	%f3, %f3, %f0
"11001100000001010000000000000001",	-- 3650: 	lli	%r5, 1
"10000100011001010010100000000000",	-- 3651: 	add	%r5, %r3, %r5
"10010000101001000000000000000000",	-- 3652: 	lf	%f4, [%r5 + 0]
"11101000011001000001100000000000",	-- 3653: 	mulf	%f3, %f3, %f4
"11001100000001010000000000000001",	-- 3654: 	lli	%r5, 1
"10000100010001010010100000000000",	-- 3655: 	add	%r5, %r2, %r5
"10010000101001000000000000000000",	-- 3656: 	lf	%f4, [%r5 + 0]
"11101000011001000010000000000000",	-- 3657: 	mulf	%f4, %f3, %f4
"11100000100000010010000000000000",	-- 3658: 	addf	%f4, %f4, %f1
"00111100100111100000000000000000",	-- 3659: 	sw	%r4, [%sp + 0]
"10110000000111100000000000000001",	-- 3660: 	sf	%f0, [%sp + 1]
"10110000001111100000000000000010",	-- 3661: 	sf	%f1, [%sp + 2]
"00111100011111100000000000000011",	-- 3662: 	sw	%r3, [%sp + 3]
"10110000010111100000000000000100",	-- 3663: 	sf	%f2, [%sp + 4]
"10110000011111100000000000000101",	-- 3664: 	sf	%f3, [%sp + 5]
"00111100010111100000000000000110",	-- 3665: 	sw	%r2, [%sp + 6]
"00111100001111100000000000000111",	-- 3666: 	sw	%r1, [%sp + 7]
"00001100100000000000000000000000",	-- 3667: 	movf	%f0, %f4
"00111111111111100000000000001000",	-- 3668: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 3669: 	addi	%sp, %sp, 9
"01011000000000000010101001001101",	-- 3670: 	jal	yj_fabs
"10101011110111100000000000001001",	-- 3671: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 3672: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000111",	-- 3673: 	lw	%r1, [%sp + 7]
"10110000000111100000000000001000",	-- 3674: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 3675: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 3676: 	addi	%sp, %sp, 10
"01011000000000000000011001011101",	-- 3677: 	jal	o_param_b.2634
"10101011110111100000000000001010",	-- 3678: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 3679: 	lw	%ra, [%sp + 9]
"00001100000000010000000000000000",	-- 3680: 	movf	%f1, %f0
"10010011110000000000000000001000",	-- 3681: 	lf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 3682: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 3683: 	addi	%sp, %sp, 10
"01011000000000000000010011110001",	-- 3684: 	jal	fless.2532
"10101011110111100000000000001010",	-- 3685: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 3686: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000000",	-- 3687: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3688: 	bneq	%r1, %r2, bneq_else.9006
"11001100000000010000000000000000",	-- 3689: 	lli	%r1, 0
"01010100000000000000111010011000",	-- 3690: 	j	bneq_cont.9007
	-- bneq_else.9006:
"11001100000000010000000000000010",	-- 3691: 	lli	%r1, 2
"00111011110000100000000000000110",	-- 3692: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 3693: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3694: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000000101",	-- 3695: 	lf	%f1, [%sp + 5]
"11101000001000000000000000000000",	-- 3696: 	mulf	%f0, %f1, %f0
"10010011110000100000000000000100",	-- 3697: 	lf	%f2, [%sp + 4]
"11100000000000100000000000000000",	-- 3698: 	addf	%f0, %f0, %f2
"00111111111111100000000000001001",	-- 3699: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 3700: 	addi	%sp, %sp, 10
"01011000000000000010101001001101",	-- 3701: 	jal	yj_fabs
"10101011110111100000000000001010",	-- 3702: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 3703: 	lw	%ra, [%sp + 9]
"00111011110000010000000000000111",	-- 3704: 	lw	%r1, [%sp + 7]
"10110000000111100000000000001001",	-- 3705: 	sf	%f0, [%sp + 9]
"00111111111111100000000000001010",	-- 3706: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 3707: 	addi	%sp, %sp, 11
"01011000000000000000011001100010",	-- 3708: 	jal	o_param_c.2636
"10101011110111100000000000001011",	-- 3709: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 3710: 	lw	%ra, [%sp + 10]
"00001100000000010000000000000000",	-- 3711: 	movf	%f1, %f0
"10010011110000000000000000001001",	-- 3712: 	lf	%f0, [%sp + 9]
"00111111111111100000000000001010",	-- 3713: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 3714: 	addi	%sp, %sp, 11
"01011000000000000000010011110001",	-- 3715: 	jal	fless.2532
"10101011110111100000000000001011",	-- 3716: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 3717: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 3718: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3719: 	bneq	%r1, %r2, bneq_else.9008
"11001100000000010000000000000000",	-- 3720: 	lli	%r1, 0
"01010100000000000000111010011000",	-- 3721: 	j	bneq_cont.9009
	-- bneq_else.9008:
"11001100000000010000000000000001",	-- 3722: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 3723: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 3724: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3725: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000001010",	-- 3726: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 3727: 	addi	%sp, %sp, 11
"01011000000000000000010011100010",	-- 3728: 	jal	fiszero.2526
"10101011110111100000000000001011",	-- 3729: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 3730: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 3731: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3732: 	bneq	%r1, %r2, bneq_else.9010
"11001100000000010000000000000001",	-- 3733: 	lli	%r1, 1
"01010100000000000000111010011000",	-- 3734: 	j	bneq_cont.9011
	-- bneq_else.9010:
"11001100000000010000000000000000",	-- 3735: 	lli	%r1, 0
	-- bneq_cont.9011:
	-- bneq_cont.9009:
	-- bneq_cont.9007:
"11001100000000100000000000000000",	-- 3736: 	lli	%r2, 0
"00101000001000100000000011000011",	-- 3737: 	bneq	%r1, %r2, bneq_else.9012
"11001100000000010000000000000010",	-- 3738: 	lli	%r1, 2
"00111011110000100000000000000011",	-- 3739: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 3740: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3741: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000000010",	-- 3742: 	lf	%f1, [%sp + 2]
"11100100000000010000000000000000",	-- 3743: 	subf	%f0, %f0, %f1
"11001100000000010000000000000011",	-- 3744: 	lli	%r1, 3
"10000100010000010000100000000000",	-- 3745: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 3746: 	lf	%f2, [%r1 + 0]
"11101000000000100000000000000000",	-- 3747: 	mulf	%f0, %f0, %f2
"11001100000000010000000000000000",	-- 3748: 	lli	%r1, 0
"00111011110000110000000000000110",	-- 3749: 	lw	%r3, [%sp + 6]
"10000100011000010000100000000000",	-- 3750: 	add	%r1, %r3, %r1
"10010000001000100000000000000000",	-- 3751: 	lf	%f2, [%r1 + 0]
"11101000000000100001000000000000",	-- 3752: 	mulf	%f2, %f0, %f2
"10010011110000110000000000000001",	-- 3753: 	lf	%f3, [%sp + 1]
"11100000010000110001000000000000",	-- 3754: 	addf	%f2, %f2, %f3
"10110000000111100000000000001010",	-- 3755: 	sf	%f0, [%sp + 10]
"00001100010000000000000000000000",	-- 3756: 	movf	%f0, %f2
"00111111111111100000000000001011",	-- 3757: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 3758: 	addi	%sp, %sp, 12
"01011000000000000010101001001101",	-- 3759: 	jal	yj_fabs
"10101011110111100000000000001100",	-- 3760: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3761: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000111",	-- 3762: 	lw	%r1, [%sp + 7]
"10110000000111100000000000001011",	-- 3763: 	sf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 3764: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3765: 	addi	%sp, %sp, 13
"01011000000000000000011001011000",	-- 3766: 	jal	o_param_a.2632
"10101011110111100000000000001101",	-- 3767: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3768: 	lw	%ra, [%sp + 12]
"00001100000000010000000000000000",	-- 3769: 	movf	%f1, %f0
"10010011110000000000000000001011",	-- 3770: 	lf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 3771: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3772: 	addi	%sp, %sp, 13
"01011000000000000000010011110001",	-- 3773: 	jal	fless.2532
"10101011110111100000000000001101",	-- 3774: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3775: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000000",	-- 3776: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3777: 	bneq	%r1, %r2, bneq_else.9013
"11001100000000010000000000000000",	-- 3778: 	lli	%r1, 0
"01010100000000000000111011110001",	-- 3779: 	j	bneq_cont.9014
	-- bneq_else.9013:
"11001100000000010000000000000010",	-- 3780: 	lli	%r1, 2
"00111011110000100000000000000110",	-- 3781: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 3782: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3783: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000001010",	-- 3784: 	lf	%f1, [%sp + 10]
"11101000001000000000000000000000",	-- 3785: 	mulf	%f0, %f1, %f0
"10010011110000100000000000000100",	-- 3786: 	lf	%f2, [%sp + 4]
"11100000000000100000000000000000",	-- 3787: 	addf	%f0, %f0, %f2
"00111111111111100000000000001100",	-- 3788: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3789: 	addi	%sp, %sp, 13
"01011000000000000010101001001101",	-- 3790: 	jal	yj_fabs
"10101011110111100000000000001101",	-- 3791: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3792: 	lw	%ra, [%sp + 12]
"00111011110000010000000000000111",	-- 3793: 	lw	%r1, [%sp + 7]
"10110000000111100000000000001100",	-- 3794: 	sf	%f0, [%sp + 12]
"00111111111111100000000000001101",	-- 3795: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 3796: 	addi	%sp, %sp, 14
"01011000000000000000011001100010",	-- 3797: 	jal	o_param_c.2636
"10101011110111100000000000001110",	-- 3798: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 3799: 	lw	%ra, [%sp + 13]
"00001100000000010000000000000000",	-- 3800: 	movf	%f1, %f0
"10010011110000000000000000001100",	-- 3801: 	lf	%f0, [%sp + 12]
"00111111111111100000000000001101",	-- 3802: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 3803: 	addi	%sp, %sp, 14
"01011000000000000000010011110001",	-- 3804: 	jal	fless.2532
"10101011110111100000000000001110",	-- 3805: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 3806: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 3807: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3808: 	bneq	%r1, %r2, bneq_else.9015
"11001100000000010000000000000000",	-- 3809: 	lli	%r1, 0
"01010100000000000000111011110001",	-- 3810: 	j	bneq_cont.9016
	-- bneq_else.9015:
"11001100000000010000000000000011",	-- 3811: 	lli	%r1, 3
"00111011110000100000000000000011",	-- 3812: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 3813: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3814: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000001101",	-- 3815: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 3816: 	addi	%sp, %sp, 14
"01011000000000000000010011100010",	-- 3817: 	jal	fiszero.2526
"10101011110111100000000000001110",	-- 3818: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 3819: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 3820: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3821: 	bneq	%r1, %r2, bneq_else.9017
"11001100000000010000000000000001",	-- 3822: 	lli	%r1, 1
"01010100000000000000111011110001",	-- 3823: 	j	bneq_cont.9018
	-- bneq_else.9017:
"11001100000000010000000000000000",	-- 3824: 	lli	%r1, 0
	-- bneq_cont.9018:
	-- bneq_cont.9016:
	-- bneq_cont.9014:
"11001100000000100000000000000000",	-- 3825: 	lli	%r2, 0
"00101000001000100000000001100011",	-- 3826: 	bneq	%r1, %r2, bneq_else.9019
"11001100000000010000000000000100",	-- 3827: 	lli	%r1, 4
"00111011110000100000000000000011",	-- 3828: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 3829: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3830: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000000100",	-- 3831: 	lf	%f1, [%sp + 4]
"11100100000000010000000000000000",	-- 3832: 	subf	%f0, %f0, %f1
"11001100000000010000000000000101",	-- 3833: 	lli	%r1, 5
"10000100010000010000100000000000",	-- 3834: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3835: 	lf	%f1, [%r1 + 0]
"11101000000000010000000000000000",	-- 3836: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000000",	-- 3837: 	lli	%r1, 0
"00111011110000110000000000000110",	-- 3838: 	lw	%r3, [%sp + 6]
"10000100011000010000100000000000",	-- 3839: 	add	%r1, %r3, %r1
"10010000001000010000000000000000",	-- 3840: 	lf	%f1, [%r1 + 0]
"11101000000000010000100000000000",	-- 3841: 	mulf	%f1, %f0, %f1
"10010011110000100000000000000001",	-- 3842: 	lf	%f2, [%sp + 1]
"11100000001000100000100000000000",	-- 3843: 	addf	%f1, %f1, %f2
"10110000000111100000000000001101",	-- 3844: 	sf	%f0, [%sp + 13]
"00001100001000000000000000000000",	-- 3845: 	movf	%f0, %f1
"00111111111111100000000000001110",	-- 3846: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 3847: 	addi	%sp, %sp, 15
"01011000000000000010101001001101",	-- 3848: 	jal	yj_fabs
"10101011110111100000000000001111",	-- 3849: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 3850: 	lw	%ra, [%sp + 14]
"00111011110000010000000000000111",	-- 3851: 	lw	%r1, [%sp + 7]
"10110000000111100000000000001110",	-- 3852: 	sf	%f0, [%sp + 14]
"00111111111111100000000000001111",	-- 3853: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 3854: 	addi	%sp, %sp, 16
"01011000000000000000011001011000",	-- 3855: 	jal	o_param_a.2632
"10101011110111100000000000010000",	-- 3856: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 3857: 	lw	%ra, [%sp + 15]
"00001100000000010000000000000000",	-- 3858: 	movf	%f1, %f0
"10010011110000000000000000001110",	-- 3859: 	lf	%f0, [%sp + 14]
"00111111111111100000000000001111",	-- 3860: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 3861: 	addi	%sp, %sp, 16
"01011000000000000000010011110001",	-- 3862: 	jal	fless.2532
"10101011110111100000000000010000",	-- 3863: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 3864: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 3865: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3866: 	bneq	%r1, %r2, bneq_else.9020
"11001100000000010000000000000000",	-- 3867: 	lli	%r1, 0
"01010100000000000000111101001010",	-- 3868: 	j	bneq_cont.9021
	-- bneq_else.9020:
"11001100000000010000000000000001",	-- 3869: 	lli	%r1, 1
"00111011110000100000000000000110",	-- 3870: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 3871: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3872: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000001101",	-- 3873: 	lf	%f1, [%sp + 13]
"11101000001000000000000000000000",	-- 3874: 	mulf	%f0, %f1, %f0
"10010011110000100000000000000010",	-- 3875: 	lf	%f2, [%sp + 2]
"11100000000000100000000000000000",	-- 3876: 	addf	%f0, %f0, %f2
"00111111111111100000000000001111",	-- 3877: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 3878: 	addi	%sp, %sp, 16
"01011000000000000010101001001101",	-- 3879: 	jal	yj_fabs
"10101011110111100000000000010000",	-- 3880: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 3881: 	lw	%ra, [%sp + 15]
"00111011110000010000000000000111",	-- 3882: 	lw	%r1, [%sp + 7]
"10110000000111100000000000001111",	-- 3883: 	sf	%f0, [%sp + 15]
"00111111111111100000000000010000",	-- 3884: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 3885: 	addi	%sp, %sp, 17
"01011000000000000000011001011101",	-- 3886: 	jal	o_param_b.2634
"10101011110111100000000000010001",	-- 3887: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 3888: 	lw	%ra, [%sp + 16]
"00001100000000010000000000000000",	-- 3889: 	movf	%f1, %f0
"10010011110000000000000000001111",	-- 3890: 	lf	%f0, [%sp + 15]
"00111111111111100000000000010000",	-- 3891: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 3892: 	addi	%sp, %sp, 17
"01011000000000000000010011110001",	-- 3893: 	jal	fless.2532
"10101011110111100000000000010001",	-- 3894: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 3895: 	lw	%ra, [%sp + 16]
"11001100000000100000000000000000",	-- 3896: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3897: 	bneq	%r1, %r2, bneq_else.9022
"11001100000000010000000000000000",	-- 3898: 	lli	%r1, 0
"01010100000000000000111101001010",	-- 3899: 	j	bneq_cont.9023
	-- bneq_else.9022:
"11001100000000010000000000000101",	-- 3900: 	lli	%r1, 5
"00111011110000100000000000000011",	-- 3901: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 3902: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3903: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000010000",	-- 3904: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 3905: 	addi	%sp, %sp, 17
"01011000000000000000010011100010",	-- 3906: 	jal	fiszero.2526
"10101011110111100000000000010001",	-- 3907: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 3908: 	lw	%ra, [%sp + 16]
"11001100000000100000000000000000",	-- 3909: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3910: 	bneq	%r1, %r2, bneq_else.9024
"11001100000000010000000000000001",	-- 3911: 	lli	%r1, 1
"01010100000000000000111101001010",	-- 3912: 	j	bneq_cont.9025
	-- bneq_else.9024:
"11001100000000010000000000000000",	-- 3913: 	lli	%r1, 0
	-- bneq_cont.9025:
	-- bneq_cont.9023:
	-- bneq_cont.9021:
"11001100000000100000000000000000",	-- 3914: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3915: 	bneq	%r1, %r2, bneq_else.9026
"11001100000000010000000000000000",	-- 3916: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3917: 	jr	%ra
	-- bneq_else.9026:
"11001100000000010000000000000000",	-- 3918: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 3919: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3920: 	add	%r1, %r2, %r1
"10010011110000000000000000001101",	-- 3921: 	lf	%f0, [%sp + 13]
"10110000000000010000000000000000",	-- 3922: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 3923: 	lli	%r1, 3
"01001111111000000000000000000000",	-- 3924: 	jr	%ra
	-- bneq_else.9019:
"11001100000000010000000000000000",	-- 3925: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 3926: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3927: 	add	%r1, %r2, %r1
"10010011110000000000000000001010",	-- 3928: 	lf	%f0, [%sp + 10]
"10110000000000010000000000000000",	-- 3929: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 3930: 	lli	%r1, 2
"01001111111000000000000000000000",	-- 3931: 	jr	%ra
	-- bneq_else.9012:
"11001100000000010000000000000000",	-- 3932: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 3933: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3934: 	add	%r1, %r2, %r1
"10010011110000000000000000000101",	-- 3935: 	lf	%f0, [%sp + 5]
"10110000000000010000000000000000",	-- 3936: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 3937: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 3938: 	jr	%ra
	-- solver_surface_fast.2767:
"00111011011000010000000000000001",	-- 3939: 	lw	%r1, [%r27 + 1]
"11001100000000110000000000000000",	-- 3940: 	lli	%r3, 0
"10000100010000110001100000000000",	-- 3941: 	add	%r3, %r2, %r3
"10010000011000110000000000000000",	-- 3942: 	lf	%f3, [%r3 + 0]
"00111100001111100000000000000000",	-- 3943: 	sw	%r1, [%sp + 0]
"10110000010111100000000000000001",	-- 3944: 	sf	%f2, [%sp + 1]
"10110000001111100000000000000010",	-- 3945: 	sf	%f1, [%sp + 2]
"10110000000111100000000000000011",	-- 3946: 	sf	%f0, [%sp + 3]
"00111100010111100000000000000100",	-- 3947: 	sw	%r2, [%sp + 4]
"00001100011000000000000000000000",	-- 3948: 	movf	%f0, %f3
"00111111111111100000000000000101",	-- 3949: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 3950: 	addi	%sp, %sp, 6
"01011000000000000000010011011011",	-- 3951: 	jal	fisneg.2524
"10101011110111100000000000000110",	-- 3952: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 3953: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000000",	-- 3954: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3955: 	bneq	%r1, %r2, bneq_else.9027
"11001100000000010000000000000000",	-- 3956: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3957: 	jr	%ra
	-- bneq_else.9027:
"11001100000000010000000000000000",	-- 3958: 	lli	%r1, 0
"11001100000000100000000000000001",	-- 3959: 	lli	%r2, 1
"00111011110000110000000000000100",	-- 3960: 	lw	%r3, [%sp + 4]
"10000100011000100001000000000000",	-- 3961: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 3962: 	lf	%f0, [%r2 + 0]
"10010011110000010000000000000011",	-- 3963: 	lf	%f1, [%sp + 3]
"11101000000000010000000000000000",	-- 3964: 	mulf	%f0, %f0, %f1
"11001100000000100000000000000010",	-- 3965: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 3966: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 3967: 	lf	%f1, [%r2 + 0]
"10010011110000100000000000000010",	-- 3968: 	lf	%f2, [%sp + 2]
"11101000001000100000100000000000",	-- 3969: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 3970: 	addf	%f0, %f0, %f1
"11001100000000100000000000000011",	-- 3971: 	lli	%r2, 3
"10000100011000100001000000000000",	-- 3972: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 3973: 	lf	%f1, [%r2 + 0]
"10010011110000100000000000000001",	-- 3974: 	lf	%f2, [%sp + 1]
"11101000001000100000100000000000",	-- 3975: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 3976: 	addf	%f0, %f0, %f1
"00111011110000100000000000000000",	-- 3977: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3978: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 3979: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 3980: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 3981: 	jr	%ra
	-- solver_second_fast.2773:
"00111011011000110000000000000001",	-- 3982: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 3983: 	lli	%r4, 0
"10000100010001000010000000000000",	-- 3984: 	add	%r4, %r2, %r4
"10010000100000110000000000000000",	-- 3985: 	lf	%f3, [%r4 + 0]
"00111100011111100000000000000000",	-- 3986: 	sw	%r3, [%sp + 0]
"10110000011111100000000000000001",	-- 3987: 	sf	%f3, [%sp + 1]
"00111100001111100000000000000010",	-- 3988: 	sw	%r1, [%sp + 2]
"10110000010111100000000000000011",	-- 3989: 	sf	%f2, [%sp + 3]
"10110000001111100000000000000100",	-- 3990: 	sf	%f1, [%sp + 4]
"10110000000111100000000000000101",	-- 3991: 	sf	%f0, [%sp + 5]
"00111100010111100000000000000110",	-- 3992: 	sw	%r2, [%sp + 6]
"00001100011000000000000000000000",	-- 3993: 	movf	%f0, %f3
"00111111111111100000000000000111",	-- 3994: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 3995: 	addi	%sp, %sp, 8
"01011000000000000000010011100010",	-- 3996: 	jal	fiszero.2526
"10101011110111100000000000001000",	-- 3997: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 3998: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000000",	-- 3999: 	lli	%r2, 0
"00101000001000100000000001110011",	-- 4000: 	bneq	%r1, %r2, bneq_else.9028
"11001100000000010000000000000001",	-- 4001: 	lli	%r1, 1
"00111011110000100000000000000110",	-- 4002: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 4003: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 4004: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000000101",	-- 4005: 	lf	%f1, [%sp + 5]
"11101000000000010000000000000000",	-- 4006: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000010",	-- 4007: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 4008: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 4009: 	lf	%f2, [%r1 + 0]
"10010011110000110000000000000100",	-- 4010: 	lf	%f3, [%sp + 4]
"11101000010000110001000000000000",	-- 4011: 	mulf	%f2, %f2, %f3
"11100000000000100000000000000000",	-- 4012: 	addf	%f0, %f0, %f2
"11001100000000010000000000000011",	-- 4013: 	lli	%r1, 3
"10000100010000010000100000000000",	-- 4014: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 4015: 	lf	%f2, [%r1 + 0]
"10010011110001000000000000000011",	-- 4016: 	lf	%f4, [%sp + 3]
"11101000010001000001000000000000",	-- 4017: 	mulf	%f2, %f2, %f4
"11100000000000100000000000000000",	-- 4018: 	addf	%f0, %f0, %f2
"00111011110000010000000000000010",	-- 4019: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000111",	-- 4020: 	sf	%f0, [%sp + 7]
"00001100100000100000000000000000",	-- 4021: 	movf	%f2, %f4
"00001100001000000000000000000000",	-- 4022: 	movf	%f0, %f1
"00001100011000010000000000000000",	-- 4023: 	movf	%f1, %f3
"00111111111111100000000000001000",	-- 4024: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 4025: 	addi	%sp, %sp, 9
"01011000000000000000110001111000",	-- 4026: 	jal	quadratic.2737
"10101011110111100000000000001001",	-- 4027: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 4028: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000010",	-- 4029: 	lw	%r1, [%sp + 2]
"10110000000111100000000000001000",	-- 4030: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 4031: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4032: 	addi	%sp, %sp, 10
"01011000000000000000011001010000",	-- 4033: 	jal	o_form.2624
"10101011110111100000000000001010",	-- 4034: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4035: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000011",	-- 4036: 	lli	%r2, 3
"00101000001000100000000000000110",	-- 4037: 	bneq	%r1, %r2, bneq_else.9029
"00010100000000000000000000000000",	-- 4038: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 4039: 	lhif	%f0, 1.000000
"10010011110000010000000000001000",	-- 4040: 	lf	%f1, [%sp + 8]
"11100100001000000000000000000000",	-- 4041: 	subf	%f0, %f1, %f0
"01010100000000000000111111001100",	-- 4042: 	j	bneq_cont.9030
	-- bneq_else.9029:
"10010011110000000000000000001000",	-- 4043: 	lf	%f0, [%sp + 8]
	-- bneq_cont.9030:
"10010011110000010000000000000111",	-- 4044: 	lf	%f1, [%sp + 7]
"10110000000111100000000000001001",	-- 4045: 	sf	%f0, [%sp + 9]
"00001100001000000000000000000000",	-- 4046: 	movf	%f0, %f1
"00111111111111100000000000001010",	-- 4047: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4048: 	addi	%sp, %sp, 11
"01011000000000000000010011101111",	-- 4049: 	jal	fsqr.2530
"10101011110111100000000000001011",	-- 4050: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4051: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 4052: 	lf	%f1, [%sp + 9]
"10010011110000100000000000000001",	-- 4053: 	lf	%f2, [%sp + 1]
"11101000010000010000100000000000",	-- 4054: 	mulf	%f1, %f2, %f1
"11100100000000010000000000000000",	-- 4055: 	subf	%f0, %f0, %f1
"10110000000111100000000000001010",	-- 4056: 	sf	%f0, [%sp + 10]
"00111111111111100000000000001011",	-- 4057: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4058: 	addi	%sp, %sp, 12
"01011000000000000000010011010100",	-- 4059: 	jal	fispos.2522
"10101011110111100000000000001100",	-- 4060: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4061: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 4062: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 4063: 	bneq	%r1, %r2, bneq_else.9031
"11001100000000010000000000000000",	-- 4064: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 4065: 	jr	%ra
	-- bneq_else.9031:
"00111011110000010000000000000010",	-- 4066: 	lw	%r1, [%sp + 2]
"00111111111111100000000000001011",	-- 4067: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4068: 	addi	%sp, %sp, 12
"01011000000000000000011001010100",	-- 4069: 	jal	o_isinvert.2628
"10101011110111100000000000001100",	-- 4070: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4071: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 4072: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 4073: 	bneq	%r1, %r2, bneq_else.9032
"11001100000000010000000000000000",	-- 4074: 	lli	%r1, 0
"10010011110000000000000000001010",	-- 4075: 	lf	%f0, [%sp + 10]
"00111100001111100000000000001011",	-- 4076: 	sw	%r1, [%sp + 11]
"00111111111111100000000000001100",	-- 4077: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4078: 	addi	%sp, %sp, 13
"01011000000000000010101000101110",	-- 4079: 	jal	yj_sqrt
"10101011110111100000000000001101",	-- 4080: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4081: 	lw	%ra, [%sp + 12]
"10010011110000010000000000000111",	-- 4082: 	lf	%f1, [%sp + 7]
"11100100001000000000000000000000",	-- 4083: 	subf	%f0, %f1, %f0
"11001100000000010000000000000100",	-- 4084: 	lli	%r1, 4
"00111011110000100000000000000110",	-- 4085: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 4086: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4087: 	lf	%f1, [%r1 + 0]
"11101000000000010000000000000000",	-- 4088: 	mulf	%f0, %f0, %f1
"00111011110000010000000000001011",	-- 4089: 	lw	%r1, [%sp + 11]
"00111011110000100000000000000000",	-- 4090: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 4091: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4092: 	sf	%f0, [%r1 + 0]
"01010100000000000001000000010001",	-- 4093: 	j	bneq_cont.9033
	-- bneq_else.9032:
"11001100000000010000000000000000",	-- 4094: 	lli	%r1, 0
"10010011110000000000000000001010",	-- 4095: 	lf	%f0, [%sp + 10]
"00111100001111100000000000001100",	-- 4096: 	sw	%r1, [%sp + 12]
"00111111111111100000000000001101",	-- 4097: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 4098: 	addi	%sp, %sp, 14
"01011000000000000010101000101110",	-- 4099: 	jal	yj_sqrt
"10101011110111100000000000001110",	-- 4100: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 4101: 	lw	%ra, [%sp + 13]
"10010011110000010000000000000111",	-- 4102: 	lf	%f1, [%sp + 7]
"11100000001000000000000000000000",	-- 4103: 	addf	%f0, %f1, %f0
"11001100000000010000000000000100",	-- 4104: 	lli	%r1, 4
"00111011110000100000000000000110",	-- 4105: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 4106: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4107: 	lf	%f1, [%r1 + 0]
"11101000000000010000000000000000",	-- 4108: 	mulf	%f0, %f0, %f1
"00111011110000010000000000001100",	-- 4109: 	lw	%r1, [%sp + 12]
"00111011110000100000000000000000",	-- 4110: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 4111: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4112: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9033:
"11001100000000010000000000000001",	-- 4113: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 4114: 	jr	%ra
	-- bneq_else.9028:
"11001100000000010000000000000000",	-- 4115: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 4116: 	jr	%ra
	-- solver_fast.2779:
"00111011011001000000000000000100",	-- 4117: 	lw	%r4, [%r27 + 4]
"00111011011001010000000000000011",	-- 4118: 	lw	%r5, [%r27 + 3]
"00111011011001100000000000000010",	-- 4119: 	lw	%r6, [%r27 + 2]
"00111011011001110000000000000001",	-- 4120: 	lw	%r7, [%r27 + 1]
"10000100111000010011100000000000",	-- 4121: 	add	%r7, %r7, %r1
"00111000111001110000000000000000",	-- 4122: 	lw	%r7, [%r7 + 0]
"11001100000010000000000000000000",	-- 4123: 	lli	%r8, 0
"10000100011010000100000000000000",	-- 4124: 	add	%r8, %r3, %r8
"10010001000000000000000000000000",	-- 4125: 	lf	%f0, [%r8 + 0]
"00111100101111100000000000000000",	-- 4126: 	sw	%r5, [%sp + 0]
"00111100100111100000000000000001",	-- 4127: 	sw	%r4, [%sp + 1]
"00111100110111100000000000000010",	-- 4128: 	sw	%r6, [%sp + 2]
"00111100001111100000000000000011",	-- 4129: 	sw	%r1, [%sp + 3]
"00111100010111100000000000000100",	-- 4130: 	sw	%r2, [%sp + 4]
"00111100111111100000000000000101",	-- 4131: 	sw	%r7, [%sp + 5]
"00111100011111100000000000000110",	-- 4132: 	sw	%r3, [%sp + 6]
"10110000000111100000000000000111",	-- 4133: 	sf	%f0, [%sp + 7]
"10000100000001110000100000000000",	-- 4134: 	add	%r1, %r0, %r7
"00111111111111100000000000001000",	-- 4135: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 4136: 	addi	%sp, %sp, 9
"01011000000000000000011001101001",	-- 4137: 	jal	o_param_x.2640
"10101011110111100000000000001001",	-- 4138: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 4139: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000111",	-- 4140: 	lf	%f1, [%sp + 7]
"11100100001000000000000000000000",	-- 4141: 	subf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 4142: 	lli	%r1, 1
"00111011110000100000000000000110",	-- 4143: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 4144: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4145: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000101",	-- 4146: 	lw	%r1, [%sp + 5]
"10110000000111100000000000001000",	-- 4147: 	sf	%f0, [%sp + 8]
"10110000001111100000000000001001",	-- 4148: 	sf	%f1, [%sp + 9]
"00111111111111100000000000001010",	-- 4149: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4150: 	addi	%sp, %sp, 11
"01011000000000000000011001101110",	-- 4151: 	jal	o_param_y.2642
"10101011110111100000000000001011",	-- 4152: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4153: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 4154: 	lf	%f1, [%sp + 9]
"11100100001000000000000000000000",	-- 4155: 	subf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 4156: 	lli	%r1, 2
"00111011110000100000000000000110",	-- 4157: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 4158: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4159: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000101",	-- 4160: 	lw	%r1, [%sp + 5]
"10110000000111100000000000001010",	-- 4161: 	sf	%f0, [%sp + 10]
"10110000001111100000000000001011",	-- 4162: 	sf	%f1, [%sp + 11]
"00111111111111100000000000001100",	-- 4163: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4164: 	addi	%sp, %sp, 13
"01011000000000000000011001110011",	-- 4165: 	jal	o_param_z.2644
"10101011110111100000000000001101",	-- 4166: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4167: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001011",	-- 4168: 	lf	%f1, [%sp + 11]
"11100100001000000000000000000000",	-- 4169: 	subf	%f0, %f1, %f0
"00111011110000010000000000000100",	-- 4170: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001100",	-- 4171: 	sf	%f0, [%sp + 12]
"00111111111111100000000000001101",	-- 4172: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 4173: 	addi	%sp, %sp, 14
"01011000000000000000011010111100",	-- 4174: 	jal	d_const.2685
"10101011110111100000000000001110",	-- 4175: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 4176: 	lw	%ra, [%sp + 13]
"00111011110000100000000000000011",	-- 4177: 	lw	%r2, [%sp + 3]
"10000100001000100000100000000000",	-- 4178: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 4179: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000000101",	-- 4180: 	lw	%r2, [%sp + 5]
"00111100001111100000000000001101",	-- 4181: 	sw	%r1, [%sp + 13]
"10000100000000100000100000000000",	-- 4182: 	add	%r1, %r0, %r2
"00111111111111100000000000001110",	-- 4183: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 4184: 	addi	%sp, %sp, 15
"01011000000000000000011001010000",	-- 4185: 	jal	o_form.2624
"10101011110111100000000000001111",	-- 4186: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 4187: 	lw	%ra, [%sp + 14]
"11001100000000100000000000000001",	-- 4188: 	lli	%r2, 1
"00101000001000100000000000010000",	-- 4189: 	bneq	%r1, %r2, bneq_else.9034
"00111011110000010000000000000100",	-- 4190: 	lw	%r1, [%sp + 4]
"00111111111111100000000000001110",	-- 4191: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 4192: 	addi	%sp, %sp, 15
"01011000000000000000011010111010",	-- 4193: 	jal	d_vec.2683
"10101011110111100000000000001111",	-- 4194: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 4195: 	lw	%ra, [%sp + 14]
"10000100000000010001000000000000",	-- 4196: 	add	%r2, %r0, %r1
"10010011110000000000000000001000",	-- 4197: 	lf	%f0, [%sp + 8]
"10010011110000010000000000001010",	-- 4198: 	lf	%f1, [%sp + 10]
"10010011110000100000000000001100",	-- 4199: 	lf	%f2, [%sp + 12]
"00111011110000010000000000000101",	-- 4200: 	lw	%r1, [%sp + 5]
"00111011110000110000000000001101",	-- 4201: 	lw	%r3, [%sp + 13]
"00111011110110110000000000000010",	-- 4202: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 4203: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 4204: 	jr	%r26
	-- bneq_else.9034:
"11001100000000100000000000000010",	-- 4205: 	lli	%r2, 2
"00101000001000100000000000001001",	-- 4206: 	bneq	%r1, %r2, bneq_else.9035
"10010011110000000000000000001000",	-- 4207: 	lf	%f0, [%sp + 8]
"10010011110000010000000000001010",	-- 4208: 	lf	%f1, [%sp + 10]
"10010011110000100000000000001100",	-- 4209: 	lf	%f2, [%sp + 12]
"00111011110000010000000000000101",	-- 4210: 	lw	%r1, [%sp + 5]
"00111011110000100000000000001101",	-- 4211: 	lw	%r2, [%sp + 13]
"00111011110110110000000000000001",	-- 4212: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 4213: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 4214: 	jr	%r26
	-- bneq_else.9035:
"10010011110000000000000000001000",	-- 4215: 	lf	%f0, [%sp + 8]
"10010011110000010000000000001010",	-- 4216: 	lf	%f1, [%sp + 10]
"10010011110000100000000000001100",	-- 4217: 	lf	%f2, [%sp + 12]
"00111011110000010000000000000101",	-- 4218: 	lw	%r1, [%sp + 5]
"00111011110000100000000000001101",	-- 4219: 	lw	%r2, [%sp + 13]
"00111011110110110000000000000000",	-- 4220: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 4221: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 4222: 	jr	%r26
	-- solver_surface_fast2.2783:
"00111011011000010000000000000001",	-- 4223: 	lw	%r1, [%r27 + 1]
"11001100000001000000000000000000",	-- 4224: 	lli	%r4, 0
"10000100010001000010000000000000",	-- 4225: 	add	%r4, %r2, %r4
"10010000100000000000000000000000",	-- 4226: 	lf	%f0, [%r4 + 0]
"00111100001111100000000000000000",	-- 4227: 	sw	%r1, [%sp + 0]
"00111100011111100000000000000001",	-- 4228: 	sw	%r3, [%sp + 1]
"00111100010111100000000000000010",	-- 4229: 	sw	%r2, [%sp + 2]
"00111111111111100000000000000011",	-- 4230: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 4231: 	addi	%sp, %sp, 4
"01011000000000000000010011011011",	-- 4232: 	jal	fisneg.2524
"10101011110111100000000000000100",	-- 4233: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 4234: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000000",	-- 4235: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 4236: 	bneq	%r1, %r2, bneq_else.9036
"11001100000000010000000000000000",	-- 4237: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 4238: 	jr	%ra
	-- bneq_else.9036:
"11001100000000010000000000000000",	-- 4239: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 4240: 	lli	%r2, 0
"00111011110000110000000000000010",	-- 4241: 	lw	%r3, [%sp + 2]
"10000100011000100001000000000000",	-- 4242: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4243: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000011",	-- 4244: 	lli	%r2, 3
"00111011110000110000000000000001",	-- 4245: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4246: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 4247: 	lf	%f1, [%r2 + 0]
"11101000000000010000000000000000",	-- 4248: 	mulf	%f0, %f0, %f1
"00111011110000100000000000000000",	-- 4249: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 4250: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4251: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 4252: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 4253: 	jr	%ra
	-- solver_second_fast2.2790:
"00111011011001000000000000000001",	-- 4254: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 4255: 	lli	%r5, 0
"10000100010001010010100000000000",	-- 4256: 	add	%r5, %r2, %r5
"10010000101000110000000000000000",	-- 4257: 	lf	%f3, [%r5 + 0]
"00111100100111100000000000000000",	-- 4258: 	sw	%r4, [%sp + 0]
"00111100001111100000000000000001",	-- 4259: 	sw	%r1, [%sp + 1]
"10110000011111100000000000000010",	-- 4260: 	sf	%f3, [%sp + 2]
"00111100011111100000000000000011",	-- 4261: 	sw	%r3, [%sp + 3]
"10110000010111100000000000000100",	-- 4262: 	sf	%f2, [%sp + 4]
"10110000001111100000000000000101",	-- 4263: 	sf	%f1, [%sp + 5]
"10110000000111100000000000000110",	-- 4264: 	sf	%f0, [%sp + 6]
"00111100010111100000000000000111",	-- 4265: 	sw	%r2, [%sp + 7]
"00001100011000000000000000000000",	-- 4266: 	movf	%f0, %f3
"00111111111111100000000000001000",	-- 4267: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 4268: 	addi	%sp, %sp, 9
"01011000000000000000010011100010",	-- 4269: 	jal	fiszero.2526
"10101011110111100000000000001001",	-- 4270: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 4271: 	lw	%ra, [%sp + 8]
"11001100000000100000000000000000",	-- 4272: 	lli	%r2, 0
"00101000001000100000000001011101",	-- 4273: 	bneq	%r1, %r2, bneq_else.9037
"11001100000000010000000000000001",	-- 4274: 	lli	%r1, 1
"00111011110000100000000000000111",	-- 4275: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 4276: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 4277: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000000110",	-- 4278: 	lf	%f1, [%sp + 6]
"11101000000000010000000000000000",	-- 4279: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000010",	-- 4280: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 4281: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4282: 	lf	%f1, [%r1 + 0]
"10010011110000100000000000000101",	-- 4283: 	lf	%f2, [%sp + 5]
"11101000001000100000100000000000",	-- 4284: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 4285: 	addf	%f0, %f0, %f1
"11001100000000010000000000000011",	-- 4286: 	lli	%r1, 3
"10000100010000010000100000000000",	-- 4287: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4288: 	lf	%f1, [%r1 + 0]
"10010011110000100000000000000100",	-- 4289: 	lf	%f2, [%sp + 4]
"11101000001000100000100000000000",	-- 4290: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 4291: 	addf	%f0, %f0, %f1
"11001100000000010000000000000011",	-- 4292: 	lli	%r1, 3
"00111011110000110000000000000011",	-- 4293: 	lw	%r3, [%sp + 3]
"10000100011000010000100000000000",	-- 4294: 	add	%r1, %r3, %r1
"10010000001000010000000000000000",	-- 4295: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000001000",	-- 4296: 	sf	%f0, [%sp + 8]
"10110000001111100000000000001001",	-- 4297: 	sf	%f1, [%sp + 9]
"00111111111111100000000000001010",	-- 4298: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4299: 	addi	%sp, %sp, 11
"01011000000000000000010011101111",	-- 4300: 	jal	fsqr.2530
"10101011110111100000000000001011",	-- 4301: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4302: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 4303: 	lf	%f1, [%sp + 9]
"10010011110000100000000000000010",	-- 4304: 	lf	%f2, [%sp + 2]
"11101000010000010000100000000000",	-- 4305: 	mulf	%f1, %f2, %f1
"11100100000000010000000000000000",	-- 4306: 	subf	%f0, %f0, %f1
"10110000000111100000000000001010",	-- 4307: 	sf	%f0, [%sp + 10]
"00111111111111100000000000001011",	-- 4308: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4309: 	addi	%sp, %sp, 12
"01011000000000000000010011010100",	-- 4310: 	jal	fispos.2522
"10101011110111100000000000001100",	-- 4311: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4312: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 4313: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 4314: 	bneq	%r1, %r2, bneq_else.9038
"11001100000000010000000000000000",	-- 4315: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 4316: 	jr	%ra
	-- bneq_else.9038:
"00111011110000010000000000000001",	-- 4317: 	lw	%r1, [%sp + 1]
"00111111111111100000000000001011",	-- 4318: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4319: 	addi	%sp, %sp, 12
"01011000000000000000011001010100",	-- 4320: 	jal	o_isinvert.2628
"10101011110111100000000000001100",	-- 4321: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4322: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 4323: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 4324: 	bneq	%r1, %r2, bneq_else.9039
"11001100000000010000000000000000",	-- 4325: 	lli	%r1, 0
"10010011110000000000000000001010",	-- 4326: 	lf	%f0, [%sp + 10]
"00111100001111100000000000001011",	-- 4327: 	sw	%r1, [%sp + 11]
"00111111111111100000000000001100",	-- 4328: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4329: 	addi	%sp, %sp, 13
"01011000000000000010101000101110",	-- 4330: 	jal	yj_sqrt
"10101011110111100000000000001101",	-- 4331: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4332: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001000",	-- 4333: 	lf	%f1, [%sp + 8]
"11100100001000000000000000000000",	-- 4334: 	subf	%f0, %f1, %f0
"11001100000000010000000000000100",	-- 4335: 	lli	%r1, 4
"00111011110000100000000000000111",	-- 4336: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 4337: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4338: 	lf	%f1, [%r1 + 0]
"11101000000000010000000000000000",	-- 4339: 	mulf	%f0, %f0, %f1
"00111011110000010000000000001011",	-- 4340: 	lw	%r1, [%sp + 11]
"00111011110000100000000000000000",	-- 4341: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 4342: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4343: 	sf	%f0, [%r1 + 0]
"01010100000000000001000100001100",	-- 4344: 	j	bneq_cont.9040
	-- bneq_else.9039:
"11001100000000010000000000000000",	-- 4345: 	lli	%r1, 0
"10010011110000000000000000001010",	-- 4346: 	lf	%f0, [%sp + 10]
"00111100001111100000000000001100",	-- 4347: 	sw	%r1, [%sp + 12]
"00111111111111100000000000001101",	-- 4348: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 4349: 	addi	%sp, %sp, 14
"01011000000000000010101000101110",	-- 4350: 	jal	yj_sqrt
"10101011110111100000000000001110",	-- 4351: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 4352: 	lw	%ra, [%sp + 13]
"10010011110000010000000000001000",	-- 4353: 	lf	%f1, [%sp + 8]
"11100000001000000000000000000000",	-- 4354: 	addf	%f0, %f1, %f0
"11001100000000010000000000000100",	-- 4355: 	lli	%r1, 4
"00111011110000100000000000000111",	-- 4356: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 4357: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4358: 	lf	%f1, [%r1 + 0]
"11101000000000010000000000000000",	-- 4359: 	mulf	%f0, %f0, %f1
"00111011110000010000000000001100",	-- 4360: 	lw	%r1, [%sp + 12]
"00111011110000100000000000000000",	-- 4361: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 4362: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4363: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9040:
"11001100000000010000000000000001",	-- 4364: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 4365: 	jr	%ra
	-- bneq_else.9037:
"11001100000000010000000000000000",	-- 4366: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 4367: 	jr	%ra
	-- solver_fast2.2797:
"00111011011000110000000000000100",	-- 4368: 	lw	%r3, [%r27 + 4]
"00111011011001000000000000000011",	-- 4369: 	lw	%r4, [%r27 + 3]
"00111011011001010000000000000010",	-- 4370: 	lw	%r5, [%r27 + 2]
"00111011011001100000000000000001",	-- 4371: 	lw	%r6, [%r27 + 1]
"10000100110000010011000000000000",	-- 4372: 	add	%r6, %r6, %r1
"00111000110001100000000000000000",	-- 4373: 	lw	%r6, [%r6 + 0]
"00111100100111100000000000000000",	-- 4374: 	sw	%r4, [%sp + 0]
"00111100011111100000000000000001",	-- 4375: 	sw	%r3, [%sp + 1]
"00111100101111100000000000000010",	-- 4376: 	sw	%r5, [%sp + 2]
"00111100110111100000000000000011",	-- 4377: 	sw	%r6, [%sp + 3]
"00111100001111100000000000000100",	-- 4378: 	sw	%r1, [%sp + 4]
"00111100010111100000000000000101",	-- 4379: 	sw	%r2, [%sp + 5]
"10000100000001100000100000000000",	-- 4380: 	add	%r1, %r0, %r6
"00111111111111100000000000000110",	-- 4381: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 4382: 	addi	%sp, %sp, 7
"01011000000000000000011010100000",	-- 4383: 	jal	o_param_ctbl.2662
"10101011110111100000000000000111",	-- 4384: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 4385: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 4386: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 4387: 	add	%r2, %r1, %r2
"10010000010000000000000000000000",	-- 4388: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000001",	-- 4389: 	lli	%r2, 1
"10000100001000100001000000000000",	-- 4390: 	add	%r2, %r1, %r2
"10010000010000010000000000000000",	-- 4391: 	lf	%f1, [%r2 + 0]
"11001100000000100000000000000010",	-- 4392: 	lli	%r2, 2
"10000100001000100001000000000000",	-- 4393: 	add	%r2, %r1, %r2
"10010000010000100000000000000000",	-- 4394: 	lf	%f2, [%r2 + 0]
"00111011110000100000000000000101",	-- 4395: 	lw	%r2, [%sp + 5]
"00111100001111100000000000000110",	-- 4396: 	sw	%r1, [%sp + 6]
"10110000010111100000000000000111",	-- 4397: 	sf	%f2, [%sp + 7]
"10110000001111100000000000001000",	-- 4398: 	sf	%f1, [%sp + 8]
"10110000000111100000000000001001",	-- 4399: 	sf	%f0, [%sp + 9]
"10000100000000100000100000000000",	-- 4400: 	add	%r1, %r0, %r2
"00111111111111100000000000001010",	-- 4401: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4402: 	addi	%sp, %sp, 11
"01011000000000000000011010111100",	-- 4403: 	jal	d_const.2685
"10101011110111100000000000001011",	-- 4404: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4405: 	lw	%ra, [%sp + 10]
"00111011110000100000000000000100",	-- 4406: 	lw	%r2, [%sp + 4]
"10000100001000100000100000000000",	-- 4407: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 4408: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000000011",	-- 4409: 	lw	%r2, [%sp + 3]
"00111100001111100000000000001010",	-- 4410: 	sw	%r1, [%sp + 10]
"10000100000000100000100000000000",	-- 4411: 	add	%r1, %r0, %r2
"00111111111111100000000000001011",	-- 4412: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4413: 	addi	%sp, %sp, 12
"01011000000000000000011001010000",	-- 4414: 	jal	o_form.2624
"10101011110111100000000000001100",	-- 4415: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4416: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000001",	-- 4417: 	lli	%r2, 1
"00101000001000100000000000010000",	-- 4418: 	bneq	%r1, %r2, bneq_else.9041
"00111011110000010000000000000101",	-- 4419: 	lw	%r1, [%sp + 5]
"00111111111111100000000000001011",	-- 4420: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4421: 	addi	%sp, %sp, 12
"01011000000000000000011010111010",	-- 4422: 	jal	d_vec.2683
"10101011110111100000000000001100",	-- 4423: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4424: 	lw	%ra, [%sp + 11]
"10000100000000010001000000000000",	-- 4425: 	add	%r2, %r0, %r1
"10010011110000000000000000001001",	-- 4426: 	lf	%f0, [%sp + 9]
"10010011110000010000000000001000",	-- 4427: 	lf	%f1, [%sp + 8]
"10010011110000100000000000000111",	-- 4428: 	lf	%f2, [%sp + 7]
"00111011110000010000000000000011",	-- 4429: 	lw	%r1, [%sp + 3]
"00111011110000110000000000001010",	-- 4430: 	lw	%r3, [%sp + 10]
"00111011110110110000000000000010",	-- 4431: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 4432: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 4433: 	jr	%r26
	-- bneq_else.9041:
"11001100000000100000000000000010",	-- 4434: 	lli	%r2, 2
"00101000001000100000000000001010",	-- 4435: 	bneq	%r1, %r2, bneq_else.9042
"10010011110000000000000000001001",	-- 4436: 	lf	%f0, [%sp + 9]
"10010011110000010000000000001000",	-- 4437: 	lf	%f1, [%sp + 8]
"10010011110000100000000000000111",	-- 4438: 	lf	%f2, [%sp + 7]
"00111011110000010000000000000011",	-- 4439: 	lw	%r1, [%sp + 3]
"00111011110000100000000000001010",	-- 4440: 	lw	%r2, [%sp + 10]
"00111011110000110000000000000110",	-- 4441: 	lw	%r3, [%sp + 6]
"00111011110110110000000000000001",	-- 4442: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 4443: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 4444: 	jr	%r26
	-- bneq_else.9042:
"10010011110000000000000000001001",	-- 4445: 	lf	%f0, [%sp + 9]
"10010011110000010000000000001000",	-- 4446: 	lf	%f1, [%sp + 8]
"10010011110000100000000000000111",	-- 4447: 	lf	%f2, [%sp + 7]
"00111011110000010000000000000011",	-- 4448: 	lw	%r1, [%sp + 3]
"00111011110000100000000000001010",	-- 4449: 	lw	%r2, [%sp + 10]
"00111011110000110000000000000110",	-- 4450: 	lw	%r3, [%sp + 6]
"00111011110110110000000000000000",	-- 4451: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 4452: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 4453: 	jr	%r26
	-- setup_rect_table.2800:
"11001100000000110000000000000110",	-- 4454: 	lli	%r3, 6
"00010100000000000000000000000000",	-- 4455: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4456: 	lhif	%f0, 0.000000
"00111100010111100000000000000000",	-- 4457: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 4458: 	sw	%r1, [%sp + 1]
"10000100000000110000100000000000",	-- 4459: 	add	%r1, %r0, %r3
"00111111111111100000000000000010",	-- 4460: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 4461: 	addi	%sp, %sp, 3
"01011000000000000010101000100010",	-- 4462: 	jal	yj_create_float_array
"10101011110111100000000000000011",	-- 4463: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 4464: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000000",	-- 4465: 	lli	%r2, 0
"00111011110000110000000000000001",	-- 4466: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4467: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4468: 	lf	%f0, [%r2 + 0]
"00111100001111100000000000000010",	-- 4469: 	sw	%r1, [%sp + 2]
"00111111111111100000000000000011",	-- 4470: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 4471: 	addi	%sp, %sp, 4
"01011000000000000000010011100010",	-- 4472: 	jal	fiszero.2526
"10101011110111100000000000000100",	-- 4473: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 4474: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000000",	-- 4475: 	lli	%r2, 0
"00101000001000100000000000111000",	-- 4476: 	bneq	%r1, %r2, bneq_else.9043
"11001100000000010000000000000000",	-- 4477: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 4478: 	lw	%r2, [%sp + 0]
"00111100001111100000000000000011",	-- 4479: 	sw	%r1, [%sp + 3]
"10000100000000100000100000000000",	-- 4480: 	add	%r1, %r0, %r2
"00111111111111100000000000000100",	-- 4481: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 4482: 	addi	%sp, %sp, 5
"01011000000000000000011001010100",	-- 4483: 	jal	o_isinvert.2628
"10101011110111100000000000000101",	-- 4484: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 4485: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000000",	-- 4486: 	lli	%r2, 0
"00111011110000110000000000000001",	-- 4487: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4488: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4489: 	lf	%f0, [%r2 + 0]
"00111100001111100000000000000100",	-- 4490: 	sw	%r1, [%sp + 4]
"00111111111111100000000000000101",	-- 4491: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 4492: 	addi	%sp, %sp, 6
"01011000000000000000010011011011",	-- 4493: 	jal	fisneg.2524
"10101011110111100000000000000110",	-- 4494: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 4495: 	lw	%ra, [%sp + 5]
"10000100000000010001000000000000",	-- 4496: 	add	%r2, %r0, %r1
"00111011110000010000000000000100",	-- 4497: 	lw	%r1, [%sp + 4]
"00111111111111100000000000000101",	-- 4498: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 4499: 	addi	%sp, %sp, 6
"01011000000000000000010011110110",	-- 4500: 	jal	xor.2565
"10101011110111100000000000000110",	-- 4501: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 4502: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000000",	-- 4503: 	lw	%r2, [%sp + 0]
"00111100001111100000000000000101",	-- 4504: 	sw	%r1, [%sp + 5]
"10000100000000100000100000000000",	-- 4505: 	add	%r1, %r0, %r2
"00111111111111100000000000000110",	-- 4506: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 4507: 	addi	%sp, %sp, 7
"01011000000000000000011001011000",	-- 4508: 	jal	o_param_a.2632
"10101011110111100000000000000111",	-- 4509: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 4510: 	lw	%ra, [%sp + 6]
"00111011110000010000000000000101",	-- 4511: 	lw	%r1, [%sp + 5]
"00111111111111100000000000000110",	-- 4512: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 4513: 	addi	%sp, %sp, 7
"01011000000000000000010100011001",	-- 4514: 	jal	fneg_cond.2570
"10101011110111100000000000000111",	-- 4515: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 4516: 	lw	%ra, [%sp + 6]
"00111011110000010000000000000011",	-- 4517: 	lw	%r1, [%sp + 3]
"00111011110000100000000000000010",	-- 4518: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4519: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4520: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 4521: 	lli	%r1, 1
"00010100000000000000000000000000",	-- 4522: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 4523: 	lhif	%f0, 1.000000
"11001100000000110000000000000000",	-- 4524: 	lli	%r3, 0
"00111011110001000000000000000001",	-- 4525: 	lw	%r4, [%sp + 1]
"10000100100000110001100000000000",	-- 4526: 	add	%r3, %r4, %r3
"10010000011000010000000000000000",	-- 4527: 	lf	%f1, [%r3 + 0]
"11101100000000010000000000000000",	-- 4528: 	divf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 4529: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4530: 	sf	%f0, [%r1 + 0]
"01010100000000000001000110111010",	-- 4531: 	j	bneq_cont.9044
	-- bneq_else.9043:
"11001100000000010000000000000001",	-- 4532: 	lli	%r1, 1
"00010100000000000000000000000000",	-- 4533: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4534: 	lhif	%f0, 0.000000
"00111011110000100000000000000010",	-- 4535: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4536: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4537: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9044:
"11001100000000010000000000000001",	-- 4538: 	lli	%r1, 1
"00111011110000110000000000000001",	-- 4539: 	lw	%r3, [%sp + 1]
"10000100011000010000100000000000",	-- 4540: 	add	%r1, %r3, %r1
"10010000001000000000000000000000",	-- 4541: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000000110",	-- 4542: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 4543: 	addi	%sp, %sp, 7
"01011000000000000000010011100010",	-- 4544: 	jal	fiszero.2526
"10101011110111100000000000000111",	-- 4545: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 4546: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 4547: 	lli	%r2, 0
"00101000001000100000000000111000",	-- 4548: 	bneq	%r1, %r2, bneq_else.9045
"11001100000000010000000000000010",	-- 4549: 	lli	%r1, 2
"00111011110000100000000000000000",	-- 4550: 	lw	%r2, [%sp + 0]
"00111100001111100000000000000110",	-- 4551: 	sw	%r1, [%sp + 6]
"10000100000000100000100000000000",	-- 4552: 	add	%r1, %r0, %r2
"00111111111111100000000000000111",	-- 4553: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 4554: 	addi	%sp, %sp, 8
"01011000000000000000011001010100",	-- 4555: 	jal	o_isinvert.2628
"10101011110111100000000000001000",	-- 4556: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 4557: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000001",	-- 4558: 	lli	%r2, 1
"00111011110000110000000000000001",	-- 4559: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4560: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4561: 	lf	%f0, [%r2 + 0]
"00111100001111100000000000000111",	-- 4562: 	sw	%r1, [%sp + 7]
"00111111111111100000000000001000",	-- 4563: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 4564: 	addi	%sp, %sp, 9
"01011000000000000000010011011011",	-- 4565: 	jal	fisneg.2524
"10101011110111100000000000001001",	-- 4566: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 4567: 	lw	%ra, [%sp + 8]
"10000100000000010001000000000000",	-- 4568: 	add	%r2, %r0, %r1
"00111011110000010000000000000111",	-- 4569: 	lw	%r1, [%sp + 7]
"00111111111111100000000000001000",	-- 4570: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 4571: 	addi	%sp, %sp, 9
"01011000000000000000010011110110",	-- 4572: 	jal	xor.2565
"10101011110111100000000000001001",	-- 4573: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 4574: 	lw	%ra, [%sp + 8]
"00111011110000100000000000000000",	-- 4575: 	lw	%r2, [%sp + 0]
"00111100001111100000000000001000",	-- 4576: 	sw	%r1, [%sp + 8]
"10000100000000100000100000000000",	-- 4577: 	add	%r1, %r0, %r2
"00111111111111100000000000001001",	-- 4578: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4579: 	addi	%sp, %sp, 10
"01011000000000000000011001011101",	-- 4580: 	jal	o_param_b.2634
"10101011110111100000000000001010",	-- 4581: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4582: 	lw	%ra, [%sp + 9]
"00111011110000010000000000001000",	-- 4583: 	lw	%r1, [%sp + 8]
"00111111111111100000000000001001",	-- 4584: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4585: 	addi	%sp, %sp, 10
"01011000000000000000010100011001",	-- 4586: 	jal	fneg_cond.2570
"10101011110111100000000000001010",	-- 4587: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4588: 	lw	%ra, [%sp + 9]
"00111011110000010000000000000110",	-- 4589: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000010",	-- 4590: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4591: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4592: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 4593: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 4594: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 4595: 	lhif	%f0, 1.000000
"11001100000000110000000000000001",	-- 4596: 	lli	%r3, 1
"00111011110001000000000000000001",	-- 4597: 	lw	%r4, [%sp + 1]
"10000100100000110001100000000000",	-- 4598: 	add	%r3, %r4, %r3
"10010000011000010000000000000000",	-- 4599: 	lf	%f1, [%r3 + 0]
"11101100000000010000000000000000",	-- 4600: 	divf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 4601: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4602: 	sf	%f0, [%r1 + 0]
"01010100000000000001001000000010",	-- 4603: 	j	bneq_cont.9046
	-- bneq_else.9045:
"11001100000000010000000000000011",	-- 4604: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 4605: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4606: 	lhif	%f0, 0.000000
"00111011110000100000000000000010",	-- 4607: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4608: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4609: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9046:
"11001100000000010000000000000010",	-- 4610: 	lli	%r1, 2
"00111011110000110000000000000001",	-- 4611: 	lw	%r3, [%sp + 1]
"10000100011000010000100000000000",	-- 4612: 	add	%r1, %r3, %r1
"10010000001000000000000000000000",	-- 4613: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000001001",	-- 4614: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4615: 	addi	%sp, %sp, 10
"01011000000000000000010011100010",	-- 4616: 	jal	fiszero.2526
"10101011110111100000000000001010",	-- 4617: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4618: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000000",	-- 4619: 	lli	%r2, 0
"00101000001000100000000000111000",	-- 4620: 	bneq	%r1, %r2, bneq_else.9047
"11001100000000010000000000000100",	-- 4621: 	lli	%r1, 4
"00111011110000100000000000000000",	-- 4622: 	lw	%r2, [%sp + 0]
"00111100001111100000000000001001",	-- 4623: 	sw	%r1, [%sp + 9]
"10000100000000100000100000000000",	-- 4624: 	add	%r1, %r0, %r2
"00111111111111100000000000001010",	-- 4625: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4626: 	addi	%sp, %sp, 11
"01011000000000000000011001010100",	-- 4627: 	jal	o_isinvert.2628
"10101011110111100000000000001011",	-- 4628: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4629: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000010",	-- 4630: 	lli	%r2, 2
"00111011110000110000000000000001",	-- 4631: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4632: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4633: 	lf	%f0, [%r2 + 0]
"00111100001111100000000000001010",	-- 4634: 	sw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 4635: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4636: 	addi	%sp, %sp, 12
"01011000000000000000010011011011",	-- 4637: 	jal	fisneg.2524
"10101011110111100000000000001100",	-- 4638: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4639: 	lw	%ra, [%sp + 11]
"10000100000000010001000000000000",	-- 4640: 	add	%r2, %r0, %r1
"00111011110000010000000000001010",	-- 4641: 	lw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 4642: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4643: 	addi	%sp, %sp, 12
"01011000000000000000010011110110",	-- 4644: 	jal	xor.2565
"10101011110111100000000000001100",	-- 4645: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4646: 	lw	%ra, [%sp + 11]
"00111011110000100000000000000000",	-- 4647: 	lw	%r2, [%sp + 0]
"00111100001111100000000000001011",	-- 4648: 	sw	%r1, [%sp + 11]
"10000100000000100000100000000000",	-- 4649: 	add	%r1, %r0, %r2
"00111111111111100000000000001100",	-- 4650: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4651: 	addi	%sp, %sp, 13
"01011000000000000000011001100010",	-- 4652: 	jal	o_param_c.2636
"10101011110111100000000000001101",	-- 4653: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4654: 	lw	%ra, [%sp + 12]
"00111011110000010000000000001011",	-- 4655: 	lw	%r1, [%sp + 11]
"00111111111111100000000000001100",	-- 4656: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4657: 	addi	%sp, %sp, 13
"01011000000000000000010100011001",	-- 4658: 	jal	fneg_cond.2570
"10101011110111100000000000001101",	-- 4659: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4660: 	lw	%ra, [%sp + 12]
"00111011110000010000000000001001",	-- 4661: 	lw	%r1, [%sp + 9]
"00111011110000100000000000000010",	-- 4662: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4663: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4664: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000101",	-- 4665: 	lli	%r1, 5
"00010100000000000000000000000000",	-- 4666: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 4667: 	lhif	%f0, 1.000000
"11001100000000110000000000000010",	-- 4668: 	lli	%r3, 2
"00111011110001000000000000000001",	-- 4669: 	lw	%r4, [%sp + 1]
"10000100100000110001100000000000",	-- 4670: 	add	%r3, %r4, %r3
"10010000011000010000000000000000",	-- 4671: 	lf	%f1, [%r3 + 0]
"11101100000000010000000000000000",	-- 4672: 	divf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 4673: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4674: 	sf	%f0, [%r1 + 0]
"01010100000000000001001001001010",	-- 4675: 	j	bneq_cont.9048
	-- bneq_else.9047:
"11001100000000010000000000000101",	-- 4676: 	lli	%r1, 5
"00010100000000000000000000000000",	-- 4677: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4678: 	lhif	%f0, 0.000000
"00111011110000100000000000000010",	-- 4679: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4680: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4681: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9048:
"10000100000000100000100000000000",	-- 4682: 	add	%r1, %r0, %r2
"01001111111000000000000000000000",	-- 4683: 	jr	%ra
	-- setup_surface_table.2803:
"11001100000000110000000000000100",	-- 4684: 	lli	%r3, 4
"00010100000000000000000000000000",	-- 4685: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4686: 	lhif	%f0, 0.000000
"00111100010111100000000000000000",	-- 4687: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 4688: 	sw	%r1, [%sp + 1]
"10000100000000110000100000000000",	-- 4689: 	add	%r1, %r0, %r3
"00111111111111100000000000000010",	-- 4690: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 4691: 	addi	%sp, %sp, 3
"01011000000000000010101000100010",	-- 4692: 	jal	yj_create_float_array
"10101011110111100000000000000011",	-- 4693: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 4694: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000000",	-- 4695: 	lli	%r2, 0
"00111011110000110000000000000001",	-- 4696: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4697: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4698: 	lf	%f0, [%r2 + 0]
"00111011110000100000000000000000",	-- 4699: 	lw	%r2, [%sp + 0]
"00111100001111100000000000000010",	-- 4700: 	sw	%r1, [%sp + 2]
"10110000000111100000000000000011",	-- 4701: 	sf	%f0, [%sp + 3]
"10000100000000100000100000000000",	-- 4702: 	add	%r1, %r0, %r2
"00111111111111100000000000000100",	-- 4703: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 4704: 	addi	%sp, %sp, 5
"01011000000000000000011001011000",	-- 4705: 	jal	o_param_a.2632
"10101011110111100000000000000101",	-- 4706: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 4707: 	lw	%ra, [%sp + 4]
"10010011110000010000000000000011",	-- 4708: 	lf	%f1, [%sp + 3]
"11101000001000000000000000000000",	-- 4709: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 4710: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 4711: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 4712: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4713: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4714: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000100",	-- 4715: 	sf	%f0, [%sp + 4]
"10110000001111100000000000000101",	-- 4716: 	sf	%f1, [%sp + 5]
"00111111111111100000000000000110",	-- 4717: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 4718: 	addi	%sp, %sp, 7
"01011000000000000000011001011101",	-- 4719: 	jal	o_param_b.2634
"10101011110111100000000000000111",	-- 4720: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 4721: 	lw	%ra, [%sp + 6]
"10010011110000010000000000000101",	-- 4722: 	lf	%f1, [%sp + 5]
"11101000001000000000000000000000",	-- 4723: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000100",	-- 4724: 	lf	%f1, [%sp + 4]
"11100000001000000000000000000000",	-- 4725: 	addf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 4726: 	lli	%r1, 2
"00111011110000100000000000000001",	-- 4727: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 4728: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4729: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4730: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000110",	-- 4731: 	sf	%f0, [%sp + 6]
"10110000001111100000000000000111",	-- 4732: 	sf	%f1, [%sp + 7]
"00111111111111100000000000001000",	-- 4733: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 4734: 	addi	%sp, %sp, 9
"01011000000000000000011001100010",	-- 4735: 	jal	o_param_c.2636
"10101011110111100000000000001001",	-- 4736: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 4737: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000111",	-- 4738: 	lf	%f1, [%sp + 7]
"11101000001000000000000000000000",	-- 4739: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000110",	-- 4740: 	lf	%f1, [%sp + 6]
"11100000001000000000000000000000",	-- 4741: 	addf	%f0, %f1, %f0
"10110000000111100000000000001000",	-- 4742: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 4743: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4744: 	addi	%sp, %sp, 10
"01011000000000000000010011010100",	-- 4745: 	jal	fispos.2522
"10101011110111100000000000001010",	-- 4746: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4747: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000000",	-- 4748: 	lli	%r2, 0
"00101000001000100000000000001000",	-- 4749: 	bneq	%r1, %r2, bneq_else.9049
"11001100000000010000000000000000",	-- 4750: 	lli	%r1, 0
"00010100000000000000000000000000",	-- 4751: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4752: 	lhif	%f0, 0.000000
"00111011110000100000000000000010",	-- 4753: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4754: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4755: 	sf	%f0, [%r1 + 0]
"01010100000000000001001011011001",	-- 4756: 	j	bneq_cont.9050
	-- bneq_else.9049:
"11001100000000010000000000000000",	-- 4757: 	lli	%r1, 0
"00010100000000000000000000000000",	-- 4758: 	llif	%f0, -1.000000
"00010000000000001011111110000000",	-- 4759: 	lhif	%f0, -1.000000
"10010011110000010000000000001000",	-- 4760: 	lf	%f1, [%sp + 8]
"11101100000000010000000000000000",	-- 4761: 	divf	%f0, %f0, %f1
"00111011110000100000000000000010",	-- 4762: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4763: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4764: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 4765: 	lli	%r1, 1
"00111011110000110000000000000000",	-- 4766: 	lw	%r3, [%sp + 0]
"00111100001111100000000000001001",	-- 4767: 	sw	%r1, [%sp + 9]
"10000100000000110000100000000000",	-- 4768: 	add	%r1, %r0, %r3
"00111111111111100000000000001010",	-- 4769: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4770: 	addi	%sp, %sp, 11
"01011000000000000000011001011000",	-- 4771: 	jal	o_param_a.2632
"10101011110111100000000000001011",	-- 4772: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4773: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001000",	-- 4774: 	lf	%f1, [%sp + 8]
"11101100000000010000000000000000",	-- 4775: 	divf	%f0, %f0, %f1
"00111111111111100000000000001010",	-- 4776: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4777: 	addi	%sp, %sp, 11
"01011000000000000010101001001111",	-- 4778: 	jal	yj_fneg
"10101011110111100000000000001011",	-- 4779: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4780: 	lw	%ra, [%sp + 10]
"00111011110000010000000000001001",	-- 4781: 	lw	%r1, [%sp + 9]
"00111011110000100000000000000010",	-- 4782: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4783: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4784: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 4785: 	lli	%r1, 2
"00111011110000110000000000000000",	-- 4786: 	lw	%r3, [%sp + 0]
"00111100001111100000000000001010",	-- 4787: 	sw	%r1, [%sp + 10]
"10000100000000110000100000000000",	-- 4788: 	add	%r1, %r0, %r3
"00111111111111100000000000001011",	-- 4789: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4790: 	addi	%sp, %sp, 12
"01011000000000000000011001011101",	-- 4791: 	jal	o_param_b.2634
"10101011110111100000000000001100",	-- 4792: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4793: 	lw	%ra, [%sp + 11]
"10010011110000010000000000001000",	-- 4794: 	lf	%f1, [%sp + 8]
"11101100000000010000000000000000",	-- 4795: 	divf	%f0, %f0, %f1
"00111111111111100000000000001011",	-- 4796: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4797: 	addi	%sp, %sp, 12
"01011000000000000010101001001111",	-- 4798: 	jal	yj_fneg
"10101011110111100000000000001100",	-- 4799: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4800: 	lw	%ra, [%sp + 11]
"00111011110000010000000000001010",	-- 4801: 	lw	%r1, [%sp + 10]
"00111011110000100000000000000010",	-- 4802: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4803: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4804: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 4805: 	lli	%r1, 3
"00111011110000110000000000000000",	-- 4806: 	lw	%r3, [%sp + 0]
"00111100001111100000000000001011",	-- 4807: 	sw	%r1, [%sp + 11]
"10000100000000110000100000000000",	-- 4808: 	add	%r1, %r0, %r3
"00111111111111100000000000001100",	-- 4809: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4810: 	addi	%sp, %sp, 13
"01011000000000000000011001100010",	-- 4811: 	jal	o_param_c.2636
"10101011110111100000000000001101",	-- 4812: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4813: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001000",	-- 4814: 	lf	%f1, [%sp + 8]
"11101100000000010000000000000000",	-- 4815: 	divf	%f0, %f0, %f1
"00111111111111100000000000001100",	-- 4816: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4817: 	addi	%sp, %sp, 13
"01011000000000000010101001001111",	-- 4818: 	jal	yj_fneg
"10101011110111100000000000001101",	-- 4819: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4820: 	lw	%ra, [%sp + 12]
"00111011110000010000000000001011",	-- 4821: 	lw	%r1, [%sp + 11]
"00111011110000100000000000000010",	-- 4822: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4823: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4824: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9050:
"10000100000000100000100000000000",	-- 4825: 	add	%r1, %r0, %r2
"01001111111000000000000000000000",	-- 4826: 	jr	%ra
	-- setup_second_table.2806:
"11001100000000110000000000000101",	-- 4827: 	lli	%r3, 5
"00010100000000000000000000000000",	-- 4828: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4829: 	lhif	%f0, 0.000000
"00111100010111100000000000000000",	-- 4830: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 4831: 	sw	%r1, [%sp + 1]
"10000100000000110000100000000000",	-- 4832: 	add	%r1, %r0, %r3
"00111111111111100000000000000010",	-- 4833: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 4834: 	addi	%sp, %sp, 3
"01011000000000000010101000100010",	-- 4835: 	jal	yj_create_float_array
"10101011110111100000000000000011",	-- 4836: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 4837: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000000",	-- 4838: 	lli	%r2, 0
"00111011110000110000000000000001",	-- 4839: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4840: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4841: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000001",	-- 4842: 	lli	%r2, 1
"10000100011000100001000000000000",	-- 4843: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 4844: 	lf	%f1, [%r2 + 0]
"11001100000000100000000000000010",	-- 4845: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 4846: 	add	%r2, %r3, %r2
"10010000010000100000000000000000",	-- 4847: 	lf	%f2, [%r2 + 0]
"00111011110000100000000000000000",	-- 4848: 	lw	%r2, [%sp + 0]
"00111100001111100000000000000010",	-- 4849: 	sw	%r1, [%sp + 2]
"10000100000000100000100000000000",	-- 4850: 	add	%r1, %r0, %r2
"00111111111111100000000000000011",	-- 4851: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 4852: 	addi	%sp, %sp, 4
"01011000000000000000110001111000",	-- 4853: 	jal	quadratic.2737
"10101011110111100000000000000100",	-- 4854: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 4855: 	lw	%ra, [%sp + 3]
"11001100000000010000000000000000",	-- 4856: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 4857: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 4858: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4859: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4860: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000011",	-- 4861: 	sf	%f0, [%sp + 3]
"10110000001111100000000000000100",	-- 4862: 	sf	%f1, [%sp + 4]
"00111111111111100000000000000101",	-- 4863: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 4864: 	addi	%sp, %sp, 6
"01011000000000000000011001011000",	-- 4865: 	jal	o_param_a.2632
"10101011110111100000000000000110",	-- 4866: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 4867: 	lw	%ra, [%sp + 5]
"10010011110000010000000000000100",	-- 4868: 	lf	%f1, [%sp + 4]
"11101000001000000000000000000000",	-- 4869: 	mulf	%f0, %f1, %f0
"00111111111111100000000000000101",	-- 4870: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 4871: 	addi	%sp, %sp, 6
"01011000000000000010101001001111",	-- 4872: 	jal	yj_fneg
"10101011110111100000000000000110",	-- 4873: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 4874: 	lw	%ra, [%sp + 5]
"11001100000000010000000000000001",	-- 4875: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 4876: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 4877: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4878: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4879: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000101",	-- 4880: 	sf	%f0, [%sp + 5]
"10110000001111100000000000000110",	-- 4881: 	sf	%f1, [%sp + 6]
"00111111111111100000000000000111",	-- 4882: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 4883: 	addi	%sp, %sp, 8
"01011000000000000000011001011101",	-- 4884: 	jal	o_param_b.2634
"10101011110111100000000000001000",	-- 4885: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 4886: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000110",	-- 4887: 	lf	%f1, [%sp + 6]
"11101000001000000000000000000000",	-- 4888: 	mulf	%f0, %f1, %f0
"00111111111111100000000000000111",	-- 4889: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 4890: 	addi	%sp, %sp, 8
"01011000000000000010101001001111",	-- 4891: 	jal	yj_fneg
"10101011110111100000000000001000",	-- 4892: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 4893: 	lw	%ra, [%sp + 7]
"11001100000000010000000000000010",	-- 4894: 	lli	%r1, 2
"00111011110000100000000000000001",	-- 4895: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 4896: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4897: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4898: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000111",	-- 4899: 	sf	%f0, [%sp + 7]
"10110000001111100000000000001000",	-- 4900: 	sf	%f1, [%sp + 8]
"00111111111111100000000000001001",	-- 4901: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4902: 	addi	%sp, %sp, 10
"01011000000000000000011001100010",	-- 4903: 	jal	o_param_c.2636
"10101011110111100000000000001010",	-- 4904: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4905: 	lw	%ra, [%sp + 9]
"10010011110000010000000000001000",	-- 4906: 	lf	%f1, [%sp + 8]
"11101000001000000000000000000000",	-- 4907: 	mulf	%f0, %f1, %f0
"00111111111111100000000000001001",	-- 4908: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4909: 	addi	%sp, %sp, 10
"01011000000000000010101001001111",	-- 4910: 	jal	yj_fneg
"10101011110111100000000000001010",	-- 4911: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4912: 	lw	%ra, [%sp + 9]
"11001100000000010000000000000000",	-- 4913: 	lli	%r1, 0
"00111011110000100000000000000010",	-- 4914: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4915: 	add	%r1, %r2, %r1
"10010011110000010000000000000011",	-- 4916: 	lf	%f1, [%sp + 3]
"10110000001000010000000000000000",	-- 4917: 	sf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4918: 	lw	%r1, [%sp + 0]
"10110000000111100000000000001001",	-- 4919: 	sf	%f0, [%sp + 9]
"00111111111111100000000000001010",	-- 4920: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4921: 	addi	%sp, %sp, 11
"01011000000000000000011001010110",	-- 4922: 	jal	o_isrot.2630
"10101011110111100000000000001011",	-- 4923: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4924: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 4925: 	lli	%r2, 0
"00101000001000100000000000001111",	-- 4926: 	bneq	%r1, %r2, bneq_else.9051
"11001100000000010000000000000001",	-- 4927: 	lli	%r1, 1
"00111011110000100000000000000010",	-- 4928: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4929: 	add	%r1, %r2, %r1
"10010011110000000000000000000101",	-- 4930: 	lf	%f0, [%sp + 5]
"10110000000000010000000000000000",	-- 4931: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 4932: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 4933: 	add	%r1, %r2, %r1
"10010011110000000000000000000111",	-- 4934: 	lf	%f0, [%sp + 7]
"10110000000000010000000000000000",	-- 4935: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 4936: 	lli	%r1, 3
"10000100010000010000100000000000",	-- 4937: 	add	%r1, %r2, %r1
"10010011110000000000000000001001",	-- 4938: 	lf	%f0, [%sp + 9]
"10110000000000010000000000000000",	-- 4939: 	sf	%f0, [%r1 + 0]
"01010100000000000001001111001110",	-- 4940: 	j	bneq_cont.9052
	-- bneq_else.9051:
"11001100000000010000000000000001",	-- 4941: 	lli	%r1, 1
"11001100000000100000000000000010",	-- 4942: 	lli	%r2, 2
"00111011110000110000000000000001",	-- 4943: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4944: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4945: 	lf	%f0, [%r2 + 0]
"00111011110000100000000000000000",	-- 4946: 	lw	%r2, [%sp + 0]
"00111100001111100000000000001010",	-- 4947: 	sw	%r1, [%sp + 10]
"10110000000111100000000000001011",	-- 4948: 	sf	%f0, [%sp + 11]
"10000100000000100000100000000000",	-- 4949: 	add	%r1, %r0, %r2
"00111111111111100000000000001100",	-- 4950: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4951: 	addi	%sp, %sp, 13
"01011000000000000000011010010110",	-- 4952: 	jal	o_param_r2.2658
"10101011110111100000000000001101",	-- 4953: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4954: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001011",	-- 4955: 	lf	%f1, [%sp + 11]
"11101000001000000000000000000000",	-- 4956: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 4957: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 4958: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 4959: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4960: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4961: 	lw	%r1, [%sp + 0]
"10110000000111100000000000001100",	-- 4962: 	sf	%f0, [%sp + 12]
"10110000001111100000000000001101",	-- 4963: 	sf	%f1, [%sp + 13]
"00111111111111100000000000001110",	-- 4964: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 4965: 	addi	%sp, %sp, 15
"01011000000000000000011010011011",	-- 4966: 	jal	o_param_r3.2660
"10101011110111100000000000001111",	-- 4967: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 4968: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001101",	-- 4969: 	lf	%f1, [%sp + 13]
"11101000001000000000000000000000",	-- 4970: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001100",	-- 4971: 	lf	%f1, [%sp + 12]
"11100000001000000000000000000000",	-- 4972: 	addf	%f0, %f1, %f0
"00111111111111100000000000001110",	-- 4973: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 4974: 	addi	%sp, %sp, 15
"01011000000000000000010011101011",	-- 4975: 	jal	fhalf.2528
"10101011110111100000000000001111",	-- 4976: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 4977: 	lw	%ra, [%sp + 14]
"10010011110000010000000000000101",	-- 4978: 	lf	%f1, [%sp + 5]
"11100100001000000000000000000000",	-- 4979: 	subf	%f0, %f1, %f0
"00111011110000010000000000001010",	-- 4980: 	lw	%r1, [%sp + 10]
"00111011110000100000000000000010",	-- 4981: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4982: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4983: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 4984: 	lli	%r1, 2
"11001100000000110000000000000010",	-- 4985: 	lli	%r3, 2
"00111011110001000000000000000001",	-- 4986: 	lw	%r4, [%sp + 1]
"10000100100000110001100000000000",	-- 4987: 	add	%r3, %r4, %r3
"10010000011000000000000000000000",	-- 4988: 	lf	%f0, [%r3 + 0]
"00111011110000110000000000000000",	-- 4989: 	lw	%r3, [%sp + 0]
"00111100001111100000000000001110",	-- 4990: 	sw	%r1, [%sp + 14]
"10110000000111100000000000001111",	-- 4991: 	sf	%f0, [%sp + 15]
"10000100000000110000100000000000",	-- 4992: 	add	%r1, %r0, %r3
"00111111111111100000000000010000",	-- 4993: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 4994: 	addi	%sp, %sp, 17
"01011000000000000000011010010001",	-- 4995: 	jal	o_param_r1.2656
"10101011110111100000000000010001",	-- 4996: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 4997: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001111",	-- 4998: 	lf	%f1, [%sp + 15]
"11101000001000000000000000000000",	-- 4999: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 5000: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 5001: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 5002: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 5003: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 5004: 	lw	%r1, [%sp + 0]
"10110000000111100000000000010000",	-- 5005: 	sf	%f0, [%sp + 16]
"10110000001111100000000000010001",	-- 5006: 	sf	%f1, [%sp + 17]
"00111111111111100000000000010010",	-- 5007: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 5008: 	addi	%sp, %sp, 19
"01011000000000000000011010011011",	-- 5009: 	jal	o_param_r3.2660
"10101011110111100000000000010011",	-- 5010: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 5011: 	lw	%ra, [%sp + 18]
"10010011110000010000000000010001",	-- 5012: 	lf	%f1, [%sp + 17]
"11101000001000000000000000000000",	-- 5013: 	mulf	%f0, %f1, %f0
"10010011110000010000000000010000",	-- 5014: 	lf	%f1, [%sp + 16]
"11100000001000000000000000000000",	-- 5015: 	addf	%f0, %f1, %f0
"00111111111111100000000000010010",	-- 5016: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 5017: 	addi	%sp, %sp, 19
"01011000000000000000010011101011",	-- 5018: 	jal	fhalf.2528
"10101011110111100000000000010011",	-- 5019: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 5020: 	lw	%ra, [%sp + 18]
"10010011110000010000000000000111",	-- 5021: 	lf	%f1, [%sp + 7]
"11100100001000000000000000000000",	-- 5022: 	subf	%f0, %f1, %f0
"00111011110000010000000000001110",	-- 5023: 	lw	%r1, [%sp + 14]
"00111011110000100000000000000010",	-- 5024: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 5025: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5026: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 5027: 	lli	%r1, 3
"11001100000000110000000000000001",	-- 5028: 	lli	%r3, 1
"00111011110001000000000000000001",	-- 5029: 	lw	%r4, [%sp + 1]
"10000100100000110001100000000000",	-- 5030: 	add	%r3, %r4, %r3
"10010000011000000000000000000000",	-- 5031: 	lf	%f0, [%r3 + 0]
"00111011110000110000000000000000",	-- 5032: 	lw	%r3, [%sp + 0]
"00111100001111100000000000010010",	-- 5033: 	sw	%r1, [%sp + 18]
"10110000000111100000000000010011",	-- 5034: 	sf	%f0, [%sp + 19]
"10000100000000110000100000000000",	-- 5035: 	add	%r1, %r0, %r3
"00111111111111100000000000010100",	-- 5036: 	sw	%ra, [%sp + 20]
"10100111110111100000000000010101",	-- 5037: 	addi	%sp, %sp, 21
"01011000000000000000011010010001",	-- 5038: 	jal	o_param_r1.2656
"10101011110111100000000000010101",	-- 5039: 	subi	%sp, %sp, 21
"00111011110111110000000000010100",	-- 5040: 	lw	%ra, [%sp + 20]
"10010011110000010000000000010011",	-- 5041: 	lf	%f1, [%sp + 19]
"11101000001000000000000000000000",	-- 5042: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 5043: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 5044: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 5045: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 5046: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 5047: 	lw	%r1, [%sp + 0]
"10110000000111100000000000010100",	-- 5048: 	sf	%f0, [%sp + 20]
"10110000001111100000000000010101",	-- 5049: 	sf	%f1, [%sp + 21]
"00111111111111100000000000010110",	-- 5050: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 5051: 	addi	%sp, %sp, 23
"01011000000000000000011010010110",	-- 5052: 	jal	o_param_r2.2658
"10101011110111100000000000010111",	-- 5053: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 5054: 	lw	%ra, [%sp + 22]
"10010011110000010000000000010101",	-- 5055: 	lf	%f1, [%sp + 21]
"11101000001000000000000000000000",	-- 5056: 	mulf	%f0, %f1, %f0
"10010011110000010000000000010100",	-- 5057: 	lf	%f1, [%sp + 20]
"11100000001000000000000000000000",	-- 5058: 	addf	%f0, %f1, %f0
"00111111111111100000000000010110",	-- 5059: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 5060: 	addi	%sp, %sp, 23
"01011000000000000000010011101011",	-- 5061: 	jal	fhalf.2528
"10101011110111100000000000010111",	-- 5062: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 5063: 	lw	%ra, [%sp + 22]
"10010011110000010000000000001001",	-- 5064: 	lf	%f1, [%sp + 9]
"11100100001000000000000000000000",	-- 5065: 	subf	%f0, %f1, %f0
"00111011110000010000000000010010",	-- 5066: 	lw	%r1, [%sp + 18]
"00111011110000100000000000000010",	-- 5067: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 5068: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5069: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9052:
"10010011110000000000000000000011",	-- 5070: 	lf	%f0, [%sp + 3]
"00111111111111100000000000010110",	-- 5071: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 5072: 	addi	%sp, %sp, 23
"01011000000000000000010011100010",	-- 5073: 	jal	fiszero.2526
"10101011110111100000000000010111",	-- 5074: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 5075: 	lw	%ra, [%sp + 22]
"11001100000000100000000000000000",	-- 5076: 	lli	%r2, 0
"00101000001000100000000000001010",	-- 5077: 	bneq	%r1, %r2, bneq_else.9053
"11001100000000010000000000000100",	-- 5078: 	lli	%r1, 4
"00010100000000000000000000000000",	-- 5079: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 5080: 	lhif	%f0, 1.000000
"10010011110000010000000000000011",	-- 5081: 	lf	%f1, [%sp + 3]
"11101100000000010000000000000000",	-- 5082: 	divf	%f0, %f0, %f1
"00111011110000100000000000000010",	-- 5083: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 5084: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5085: 	sf	%f0, [%r1 + 0]
"01010100000000000001001111011111",	-- 5086: 	j	bneq_cont.9054
	-- bneq_else.9053:
	-- bneq_cont.9054:
"00111011110000010000000000000010",	-- 5087: 	lw	%r1, [%sp + 2]
"01001111111000000000000000000000",	-- 5088: 	jr	%ra
	-- iter_setup_dirvec_constants.2809:
"00111011011000110000000000000001",	-- 5089: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 5090: 	lli	%r4, 0
"00110000100000100000000001001001",	-- 5091: 	bgt	%r4, %r2, bgt_else.9055
"10000100011000100001100000000000",	-- 5092: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 5093: 	lw	%r3, [%r3 + 0]
"00111111011111100000000000000000",	-- 5094: 	sw	%r27, [%sp + 0]
"00111100010111100000000000000001",	-- 5095: 	sw	%r2, [%sp + 1]
"00111100011111100000000000000010",	-- 5096: 	sw	%r3, [%sp + 2]
"00111100001111100000000000000011",	-- 5097: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 5098: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5099: 	addi	%sp, %sp, 5
"01011000000000000000011010111100",	-- 5100: 	jal	d_const.2685
"10101011110111100000000000000101",	-- 5101: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5102: 	lw	%ra, [%sp + 4]
"00111011110000100000000000000011",	-- 5103: 	lw	%r2, [%sp + 3]
"00111100001111100000000000000100",	-- 5104: 	sw	%r1, [%sp + 4]
"10000100000000100000100000000000",	-- 5105: 	add	%r1, %r0, %r2
"00111111111111100000000000000101",	-- 5106: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5107: 	addi	%sp, %sp, 6
"01011000000000000000011010111010",	-- 5108: 	jal	d_vec.2683
"10101011110111100000000000000110",	-- 5109: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5110: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000010",	-- 5111: 	lw	%r2, [%sp + 2]
"00111100001111100000000000000101",	-- 5112: 	sw	%r1, [%sp + 5]
"10000100000000100000100000000000",	-- 5113: 	add	%r1, %r0, %r2
"00111111111111100000000000000110",	-- 5114: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5115: 	addi	%sp, %sp, 7
"01011000000000000000011001010000",	-- 5116: 	jal	o_form.2624
"10101011110111100000000000000111",	-- 5117: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5118: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000001",	-- 5119: 	lli	%r2, 1
"00101000001000100000000000001101",	-- 5120: 	bneq	%r1, %r2, bneq_else.9056
"00111011110000010000000000000101",	-- 5121: 	lw	%r1, [%sp + 5]
"00111011110000100000000000000010",	-- 5122: 	lw	%r2, [%sp + 2]
"00111111111111100000000000000110",	-- 5123: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5124: 	addi	%sp, %sp, 7
"01011000000000000001000101100110",	-- 5125: 	jal	setup_rect_table.2800
"10101011110111100000000000000111",	-- 5126: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5127: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000001",	-- 5128: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000100",	-- 5129: 	lw	%r3, [%sp + 4]
"10000100011000100001100000000000",	-- 5130: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 5131: 	sw	%r1, [%r3 + 0]
"01010100000000000001010000100110",	-- 5132: 	j	bneq_cont.9057
	-- bneq_else.9056:
"11001100000000100000000000000010",	-- 5133: 	lli	%r2, 2
"00101000001000100000000000001101",	-- 5134: 	bneq	%r1, %r2, bneq_else.9058
"00111011110000010000000000000101",	-- 5135: 	lw	%r1, [%sp + 5]
"00111011110000100000000000000010",	-- 5136: 	lw	%r2, [%sp + 2]
"00111111111111100000000000000110",	-- 5137: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5138: 	addi	%sp, %sp, 7
"01011000000000000001001001001100",	-- 5139: 	jal	setup_surface_table.2803
"10101011110111100000000000000111",	-- 5140: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5141: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000001",	-- 5142: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000100",	-- 5143: 	lw	%r3, [%sp + 4]
"10000100011000100001100000000000",	-- 5144: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 5145: 	sw	%r1, [%r3 + 0]
"01010100000000000001010000100110",	-- 5146: 	j	bneq_cont.9059
	-- bneq_else.9058:
"00111011110000010000000000000101",	-- 5147: 	lw	%r1, [%sp + 5]
"00111011110000100000000000000010",	-- 5148: 	lw	%r2, [%sp + 2]
"00111111111111100000000000000110",	-- 5149: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5150: 	addi	%sp, %sp, 7
"01011000000000000001001011011011",	-- 5151: 	jal	setup_second_table.2806
"10101011110111100000000000000111",	-- 5152: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5153: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000001",	-- 5154: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000100",	-- 5155: 	lw	%r3, [%sp + 4]
"10000100011000100001100000000000",	-- 5156: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 5157: 	sw	%r1, [%r3 + 0]
	-- bneq_cont.9059:
	-- bneq_cont.9057:
"11001100000000010000000000000001",	-- 5158: 	lli	%r1, 1
"10001000010000010001000000000000",	-- 5159: 	sub	%r2, %r2, %r1
"00111011110000010000000000000011",	-- 5160: 	lw	%r1, [%sp + 3]
"00111011110110110000000000000000",	-- 5161: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 5162: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5163: 	jr	%r26
	-- bgt_else.9055:
"01001111111000000000000000000000",	-- 5164: 	jr	%ra
	-- setup_dirvec_constants.2812:
"00111011011000100000000000000010",	-- 5165: 	lw	%r2, [%r27 + 2]
"00111011011110110000000000000001",	-- 5166: 	lw	%r27, [%r27 + 1]
"11001100000000110000000000000000",	-- 5167: 	lli	%r3, 0
"10000100010000110001000000000000",	-- 5168: 	add	%r2, %r2, %r3
"00111000010000100000000000000000",	-- 5169: 	lw	%r2, [%r2 + 0]
"11001100000000110000000000000001",	-- 5170: 	lli	%r3, 1
"10001000010000110001000000000000",	-- 5171: 	sub	%r2, %r2, %r3
"00111011011110100000000000000000",	-- 5172: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5173: 	jr	%r26
	-- setup_startp_constants.2814:
"00111011011000110000000000000001",	-- 5174: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 5175: 	lli	%r4, 0
"00110000100000100000000010010110",	-- 5176: 	bgt	%r4, %r2, bgt_else.9061
"10000100011000100001100000000000",	-- 5177: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 5178: 	lw	%r3, [%r3 + 0]
"00111111011111100000000000000000",	-- 5179: 	sw	%r27, [%sp + 0]
"00111100010111100000000000000001",	-- 5180: 	sw	%r2, [%sp + 1]
"00111100001111100000000000000010",	-- 5181: 	sw	%r1, [%sp + 2]
"00111100011111100000000000000011",	-- 5182: 	sw	%r3, [%sp + 3]
"10000100000000110000100000000000",	-- 5183: 	add	%r1, %r0, %r3
"00111111111111100000000000000100",	-- 5184: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5185: 	addi	%sp, %sp, 5
"01011000000000000000011010100000",	-- 5186: 	jal	o_param_ctbl.2662
"10101011110111100000000000000101",	-- 5187: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5188: 	lw	%ra, [%sp + 4]
"00111011110000100000000000000011",	-- 5189: 	lw	%r2, [%sp + 3]
"00111100001111100000000000000100",	-- 5190: 	sw	%r1, [%sp + 4]
"10000100000000100000100000000000",	-- 5191: 	add	%r1, %r0, %r2
"00111111111111100000000000000101",	-- 5192: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5193: 	addi	%sp, %sp, 6
"01011000000000000000011001010000",	-- 5194: 	jal	o_form.2624
"10101011110111100000000000000110",	-- 5195: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5196: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000000",	-- 5197: 	lli	%r2, 0
"11001100000000110000000000000000",	-- 5198: 	lli	%r3, 0
"00111011110001000000000000000010",	-- 5199: 	lw	%r4, [%sp + 2]
"10000100100000110001100000000000",	-- 5200: 	add	%r3, %r4, %r3
"10010000011000000000000000000000",	-- 5201: 	lf	%f0, [%r3 + 0]
"00111011110000110000000000000011",	-- 5202: 	lw	%r3, [%sp + 3]
"00111100001111100000000000000101",	-- 5203: 	sw	%r1, [%sp + 5]
"00111100010111100000000000000110",	-- 5204: 	sw	%r2, [%sp + 6]
"10110000000111100000000000000111",	-- 5205: 	sf	%f0, [%sp + 7]
"10000100000000110000100000000000",	-- 5206: 	add	%r1, %r0, %r3
"00111111111111100000000000001000",	-- 5207: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 5208: 	addi	%sp, %sp, 9
"01011000000000000000011001101001",	-- 5209: 	jal	o_param_x.2640
"10101011110111100000000000001001",	-- 5210: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 5211: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000111",	-- 5212: 	lf	%f1, [%sp + 7]
"11100100001000000000000000000000",	-- 5213: 	subf	%f0, %f1, %f0
"00111011110000010000000000000110",	-- 5214: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000100",	-- 5215: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5216: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5217: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 5218: 	lli	%r1, 1
"11001100000000110000000000000001",	-- 5219: 	lli	%r3, 1
"00111011110001000000000000000010",	-- 5220: 	lw	%r4, [%sp + 2]
"10000100100000110001100000000000",	-- 5221: 	add	%r3, %r4, %r3
"10010000011000000000000000000000",	-- 5222: 	lf	%f0, [%r3 + 0]
"00111011110000110000000000000011",	-- 5223: 	lw	%r3, [%sp + 3]
"00111100001111100000000000001000",	-- 5224: 	sw	%r1, [%sp + 8]
"10110000000111100000000000001001",	-- 5225: 	sf	%f0, [%sp + 9]
"10000100000000110000100000000000",	-- 5226: 	add	%r1, %r0, %r3
"00111111111111100000000000001010",	-- 5227: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 5228: 	addi	%sp, %sp, 11
"01011000000000000000011001101110",	-- 5229: 	jal	o_param_y.2642
"10101011110111100000000000001011",	-- 5230: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 5231: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 5232: 	lf	%f1, [%sp + 9]
"11100100001000000000000000000000",	-- 5233: 	subf	%f0, %f1, %f0
"00111011110000010000000000001000",	-- 5234: 	lw	%r1, [%sp + 8]
"00111011110000100000000000000100",	-- 5235: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5236: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5237: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 5238: 	lli	%r1, 2
"11001100000000110000000000000010",	-- 5239: 	lli	%r3, 2
"00111011110001000000000000000010",	-- 5240: 	lw	%r4, [%sp + 2]
"10000100100000110001100000000000",	-- 5241: 	add	%r3, %r4, %r3
"10010000011000000000000000000000",	-- 5242: 	lf	%f0, [%r3 + 0]
"00111011110000110000000000000011",	-- 5243: 	lw	%r3, [%sp + 3]
"00111100001111100000000000001010",	-- 5244: 	sw	%r1, [%sp + 10]
"10110000000111100000000000001011",	-- 5245: 	sf	%f0, [%sp + 11]
"10000100000000110000100000000000",	-- 5246: 	add	%r1, %r0, %r3
"00111111111111100000000000001100",	-- 5247: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 5248: 	addi	%sp, %sp, 13
"01011000000000000000011001110011",	-- 5249: 	jal	o_param_z.2644
"10101011110111100000000000001101",	-- 5250: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 5251: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001011",	-- 5252: 	lf	%f1, [%sp + 11]
"11100100001000000000000000000000",	-- 5253: 	subf	%f0, %f1, %f0
"00111011110000010000000000001010",	-- 5254: 	lw	%r1, [%sp + 10]
"00111011110000100000000000000100",	-- 5255: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5256: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5257: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 5258: 	lli	%r1, 2
"00111011110000110000000000000101",	-- 5259: 	lw	%r3, [%sp + 5]
"00101000011000010000000000011110",	-- 5260: 	bneq	%r3, %r1, bneq_else.9062
"11001100000000010000000000000011",	-- 5261: 	lli	%r1, 3
"00111011110000110000000000000011",	-- 5262: 	lw	%r3, [%sp + 3]
"00111100001111100000000000001100",	-- 5263: 	sw	%r1, [%sp + 12]
"10000100000000110000100000000000",	-- 5264: 	add	%r1, %r0, %r3
"00111111111111100000000000001101",	-- 5265: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 5266: 	addi	%sp, %sp, 14
"01011000000000000000011001100111",	-- 5267: 	jal	o_param_abc.2638
"10101011110111100000000000001110",	-- 5268: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 5269: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 5270: 	lli	%r2, 0
"00111011110000110000000000000100",	-- 5271: 	lw	%r3, [%sp + 4]
"10000100011000100001000000000000",	-- 5272: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 5273: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000001",	-- 5274: 	lli	%r2, 1
"10000100011000100001000000000000",	-- 5275: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 5276: 	lf	%f1, [%r2 + 0]
"11001100000000100000000000000010",	-- 5277: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 5278: 	add	%r2, %r3, %r2
"10010000010000100000000000000000",	-- 5279: 	lf	%f2, [%r2 + 0]
"00111111111111100000000000001101",	-- 5280: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 5281: 	addi	%sp, %sp, 14
"01011000000000000000010110111101",	-- 5282: 	jal	veciprod2.2600
"10101011110111100000000000001110",	-- 5283: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 5284: 	lw	%ra, [%sp + 13]
"00111011110000010000000000001100",	-- 5285: 	lw	%r1, [%sp + 12]
"00111011110000100000000000000100",	-- 5286: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5287: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5288: 	sf	%f0, [%r1 + 0]
"01010100000000000001010011000111",	-- 5289: 	j	bneq_cont.9063
	-- bneq_else.9062:
"11001100000000010000000000000010",	-- 5290: 	lli	%r1, 2
"00110000011000010000000000000010",	-- 5291: 	bgt	%r3, %r1, bgt_else.9064
"01010100000000000001010011000111",	-- 5292: 	j	bgt_cont.9065
	-- bgt_else.9064:
"11001100000000010000000000000000",	-- 5293: 	lli	%r1, 0
"10000100010000010000100000000000",	-- 5294: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 5295: 	lf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 5296: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 5297: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 5298: 	lf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 5299: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 5300: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 5301: 	lf	%f2, [%r1 + 0]
"00111011110000010000000000000011",	-- 5302: 	lw	%r1, [%sp + 3]
"00111111111111100000000000001101",	-- 5303: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 5304: 	addi	%sp, %sp, 14
"01011000000000000000110001111000",	-- 5305: 	jal	quadratic.2737
"10101011110111100000000000001110",	-- 5306: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 5307: 	lw	%ra, [%sp + 13]
"11001100000000010000000000000011",	-- 5308: 	lli	%r1, 3
"11001100000000100000000000000011",	-- 5309: 	lli	%r2, 3
"00111011110000110000000000000101",	-- 5310: 	lw	%r3, [%sp + 5]
"00101000011000100000000000000101",	-- 5311: 	bneq	%r3, %r2, bneq_else.9066
"00010100000000010000000000000000",	-- 5312: 	llif	%f1, 1.000000
"00010000000000010011111110000000",	-- 5313: 	lhif	%f1, 1.000000
"11100100000000010000000000000000",	-- 5314: 	subf	%f0, %f0, %f1
"01010100000000000001010011000100",	-- 5315: 	j	bneq_cont.9067
	-- bneq_else.9066:
	-- bneq_cont.9067:
"00111011110000100000000000000100",	-- 5316: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5317: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5318: 	sf	%f0, [%r1 + 0]
	-- bgt_cont.9065:
	-- bneq_cont.9063:
"11001100000000010000000000000001",	-- 5319: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 5320: 	lw	%r2, [%sp + 1]
"10001000010000010001000000000000",	-- 5321: 	sub	%r2, %r2, %r1
"00111011110000010000000000000010",	-- 5322: 	lw	%r1, [%sp + 2]
"00111011110110110000000000000000",	-- 5323: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 5324: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5325: 	jr	%r26
	-- bgt_else.9061:
"01001111111000000000000000000000",	-- 5326: 	jr	%ra
	-- setup_startp.2817:
"00111011011000100000000000000011",	-- 5327: 	lw	%r2, [%r27 + 3]
"00111011011000110000000000000010",	-- 5328: 	lw	%r3, [%r27 + 2]
"00111011011001000000000000000001",	-- 5329: 	lw	%r4, [%r27 + 1]
"00111100001111100000000000000000",	-- 5330: 	sw	%r1, [%sp + 0]
"00111100011111100000000000000001",	-- 5331: 	sw	%r3, [%sp + 1]
"00111100100111100000000000000010",	-- 5332: 	sw	%r4, [%sp + 2]
"10000100000000101101000000000000",	-- 5333: 	add	%r26, %r0, %r2
"10000100000000010001000000000000",	-- 5334: 	add	%r2, %r0, %r1
"10000100000110100000100000000000",	-- 5335: 	add	%r1, %r0, %r26
"00111111111111100000000000000011",	-- 5336: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 5337: 	addi	%sp, %sp, 4
"01011000000000000000010100111011",	-- 5338: 	jal	veccpy.2586
"10101011110111100000000000000100",	-- 5339: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 5340: 	lw	%ra, [%sp + 3]
"11001100000000010000000000000000",	-- 5341: 	lli	%r1, 0
"00111011110000100000000000000010",	-- 5342: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 5343: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 5344: 	lw	%r1, [%r1 + 0]
"11001100000000100000000000000001",	-- 5345: 	lli	%r2, 1
"10001000001000100001000000000000",	-- 5346: 	sub	%r2, %r1, %r2
"00111011110000010000000000000000",	-- 5347: 	lw	%r1, [%sp + 0]
"00111011110110110000000000000001",	-- 5348: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 5349: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5350: 	jr	%r26
	-- is_rect_outside.2819:
"10110000010111100000000000000000",	-- 5351: 	sf	%f2, [%sp + 0]
"10110000001111100000000000000001",	-- 5352: 	sf	%f1, [%sp + 1]
"00111100001111100000000000000010",	-- 5353: 	sw	%r1, [%sp + 2]
"00111111111111100000000000000011",	-- 5354: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 5355: 	addi	%sp, %sp, 4
"01011000000000000010101001001101",	-- 5356: 	jal	yj_fabs
"10101011110111100000000000000100",	-- 5357: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 5358: 	lw	%ra, [%sp + 3]
"00111011110000010000000000000010",	-- 5359: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000011",	-- 5360: 	sf	%f0, [%sp + 3]
"00111111111111100000000000000100",	-- 5361: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5362: 	addi	%sp, %sp, 5
"01011000000000000000011001011000",	-- 5363: 	jal	o_param_a.2632
"10101011110111100000000000000101",	-- 5364: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5365: 	lw	%ra, [%sp + 4]
"00001100000000010000000000000000",	-- 5366: 	movf	%f1, %f0
"10010011110000000000000000000011",	-- 5367: 	lf	%f0, [%sp + 3]
"00111111111111100000000000000100",	-- 5368: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5369: 	addi	%sp, %sp, 5
"01011000000000000000010011110001",	-- 5370: 	jal	fless.2532
"10101011110111100000000000000101",	-- 5371: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5372: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000000",	-- 5373: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5374: 	bneq	%r1, %r2, bneq_else.9069
"11001100000000010000000000000000",	-- 5375: 	lli	%r1, 0
"01010100000000000001010100101101",	-- 5376: 	j	bneq_cont.9070
	-- bneq_else.9069:
"10010011110000000000000000000001",	-- 5377: 	lf	%f0, [%sp + 1]
"00111111111111100000000000000100",	-- 5378: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5379: 	addi	%sp, %sp, 5
"01011000000000000010101001001101",	-- 5380: 	jal	yj_fabs
"10101011110111100000000000000101",	-- 5381: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5382: 	lw	%ra, [%sp + 4]
"00111011110000010000000000000010",	-- 5383: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000100",	-- 5384: 	sf	%f0, [%sp + 4]
"00111111111111100000000000000101",	-- 5385: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5386: 	addi	%sp, %sp, 6
"01011000000000000000011001011101",	-- 5387: 	jal	o_param_b.2634
"10101011110111100000000000000110",	-- 5388: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5389: 	lw	%ra, [%sp + 5]
"00001100000000010000000000000000",	-- 5390: 	movf	%f1, %f0
"10010011110000000000000000000100",	-- 5391: 	lf	%f0, [%sp + 4]
"00111111111111100000000000000101",	-- 5392: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5393: 	addi	%sp, %sp, 6
"01011000000000000000010011110001",	-- 5394: 	jal	fless.2532
"10101011110111100000000000000110",	-- 5395: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5396: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000000",	-- 5397: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5398: 	bneq	%r1, %r2, bneq_else.9071
"11001100000000010000000000000000",	-- 5399: 	lli	%r1, 0
"01010100000000000001010100101101",	-- 5400: 	j	bneq_cont.9072
	-- bneq_else.9071:
"10010011110000000000000000000000",	-- 5401: 	lf	%f0, [%sp + 0]
"00111111111111100000000000000101",	-- 5402: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5403: 	addi	%sp, %sp, 6
"01011000000000000010101001001101",	-- 5404: 	jal	yj_fabs
"10101011110111100000000000000110",	-- 5405: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5406: 	lw	%ra, [%sp + 5]
"00111011110000010000000000000010",	-- 5407: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000101",	-- 5408: 	sf	%f0, [%sp + 5]
"00111111111111100000000000000110",	-- 5409: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5410: 	addi	%sp, %sp, 7
"01011000000000000000011001100010",	-- 5411: 	jal	o_param_c.2636
"10101011110111100000000000000111",	-- 5412: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5413: 	lw	%ra, [%sp + 6]
"00001100000000010000000000000000",	-- 5414: 	movf	%f1, %f0
"10010011110000000000000000000101",	-- 5415: 	lf	%f0, [%sp + 5]
"00111111111111100000000000000110",	-- 5416: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5417: 	addi	%sp, %sp, 7
"01011000000000000000010011110001",	-- 5418: 	jal	fless.2532
"10101011110111100000000000000111",	-- 5419: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5420: 	lw	%ra, [%sp + 6]
	-- bneq_cont.9072:
	-- bneq_cont.9070:
"11001100000000100000000000000000",	-- 5421: 	lli	%r2, 0
"00101000001000100000000000001101",	-- 5422: 	bneq	%r1, %r2, bneq_else.9073
"00111011110000010000000000000010",	-- 5423: 	lw	%r1, [%sp + 2]
"00111111111111100000000000000110",	-- 5424: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5425: 	addi	%sp, %sp, 7
"01011000000000000000011001010100",	-- 5426: 	jal	o_isinvert.2628
"10101011110111100000000000000111",	-- 5427: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5428: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5429: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5430: 	bneq	%r1, %r2, bneq_else.9074
"11001100000000010000000000000001",	-- 5431: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5432: 	jr	%ra
	-- bneq_else.9074:
"11001100000000010000000000000000",	-- 5433: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5434: 	jr	%ra
	-- bneq_else.9073:
"00111011110000010000000000000010",	-- 5435: 	lw	%r1, [%sp + 2]
"01010100000000000000011001010100",	-- 5436: 	j	o_isinvert.2628
	-- is_plane_outside.2824:
"00111100001111100000000000000000",	-- 5437: 	sw	%r1, [%sp + 0]
"10110000010111100000000000000001",	-- 5438: 	sf	%f2, [%sp + 1]
"10110000001111100000000000000010",	-- 5439: 	sf	%f1, [%sp + 2]
"10110000000111100000000000000011",	-- 5440: 	sf	%f0, [%sp + 3]
"00111111111111100000000000000100",	-- 5441: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5442: 	addi	%sp, %sp, 5
"01011000000000000000011001100111",	-- 5443: 	jal	o_param_abc.2638
"10101011110111100000000000000101",	-- 5444: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5445: 	lw	%ra, [%sp + 4]
"10010011110000000000000000000011",	-- 5446: 	lf	%f0, [%sp + 3]
"10010011110000010000000000000010",	-- 5447: 	lf	%f1, [%sp + 2]
"10010011110000100000000000000001",	-- 5448: 	lf	%f2, [%sp + 1]
"00111111111111100000000000000100",	-- 5449: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5450: 	addi	%sp, %sp, 5
"01011000000000000000010110111101",	-- 5451: 	jal	veciprod2.2600
"10101011110111100000000000000101",	-- 5452: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5453: 	lw	%ra, [%sp + 4]
"00111011110000010000000000000000",	-- 5454: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000100",	-- 5455: 	sf	%f0, [%sp + 4]
"00111111111111100000000000000101",	-- 5456: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5457: 	addi	%sp, %sp, 6
"01011000000000000000011001010100",	-- 5458: 	jal	o_isinvert.2628
"10101011110111100000000000000110",	-- 5459: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5460: 	lw	%ra, [%sp + 5]
"10010011110000000000000000000100",	-- 5461: 	lf	%f0, [%sp + 4]
"00111100001111100000000000000101",	-- 5462: 	sw	%r1, [%sp + 5]
"00111111111111100000000000000110",	-- 5463: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5464: 	addi	%sp, %sp, 7
"01011000000000000000010011011011",	-- 5465: 	jal	fisneg.2524
"10101011110111100000000000000111",	-- 5466: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5467: 	lw	%ra, [%sp + 6]
"10000100000000010001000000000000",	-- 5468: 	add	%r2, %r0, %r1
"00111011110000010000000000000101",	-- 5469: 	lw	%r1, [%sp + 5]
"00111111111111100000000000000110",	-- 5470: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5471: 	addi	%sp, %sp, 7
"01011000000000000000010011110110",	-- 5472: 	jal	xor.2565
"10101011110111100000000000000111",	-- 5473: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5474: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5475: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5476: 	bneq	%r1, %r2, bneq_else.9075
"11001100000000010000000000000001",	-- 5477: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5478: 	jr	%ra
	-- bneq_else.9075:
"11001100000000010000000000000000",	-- 5479: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5480: 	jr	%ra
	-- is_second_outside.2829:
"00111100001111100000000000000000",	-- 5481: 	sw	%r1, [%sp + 0]
"00111111111111100000000000000001",	-- 5482: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 5483: 	addi	%sp, %sp, 2
"01011000000000000000110001111000",	-- 5484: 	jal	quadratic.2737
"10101011110111100000000000000010",	-- 5485: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 5486: 	lw	%ra, [%sp + 1]
"00111011110000010000000000000000",	-- 5487: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000001",	-- 5488: 	sf	%f0, [%sp + 1]
"00111111111111100000000000000010",	-- 5489: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 5490: 	addi	%sp, %sp, 3
"01011000000000000000011001010000",	-- 5491: 	jal	o_form.2624
"10101011110111100000000000000011",	-- 5492: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 5493: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000011",	-- 5494: 	lli	%r2, 3
"00101000001000100000000000000110",	-- 5495: 	bneq	%r1, %r2, bneq_else.9076
"00010100000000000000000000000000",	-- 5496: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 5497: 	lhif	%f0, 1.000000
"10010011110000010000000000000001",	-- 5498: 	lf	%f1, [%sp + 1]
"11100100001000000000000000000000",	-- 5499: 	subf	%f0, %f1, %f0
"01010100000000000001010101111110",	-- 5500: 	j	bneq_cont.9077
	-- bneq_else.9076:
"10010011110000000000000000000001",	-- 5501: 	lf	%f0, [%sp + 1]
	-- bneq_cont.9077:
"00111011110000010000000000000000",	-- 5502: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000010",	-- 5503: 	sf	%f0, [%sp + 2]
"00111111111111100000000000000011",	-- 5504: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 5505: 	addi	%sp, %sp, 4
"01011000000000000000011001010100",	-- 5506: 	jal	o_isinvert.2628
"10101011110111100000000000000100",	-- 5507: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 5508: 	lw	%ra, [%sp + 3]
"10010011110000000000000000000010",	-- 5509: 	lf	%f0, [%sp + 2]
"00111100001111100000000000000011",	-- 5510: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 5511: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5512: 	addi	%sp, %sp, 5
"01011000000000000000010011011011",	-- 5513: 	jal	fisneg.2524
"10101011110111100000000000000101",	-- 5514: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5515: 	lw	%ra, [%sp + 4]
"10000100000000010001000000000000",	-- 5516: 	add	%r2, %r0, %r1
"00111011110000010000000000000011",	-- 5517: 	lw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 5518: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5519: 	addi	%sp, %sp, 5
"01011000000000000000010011110110",	-- 5520: 	jal	xor.2565
"10101011110111100000000000000101",	-- 5521: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5522: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000000",	-- 5523: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5524: 	bneq	%r1, %r2, bneq_else.9078
"11001100000000010000000000000001",	-- 5525: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5526: 	jr	%ra
	-- bneq_else.9078:
"11001100000000010000000000000000",	-- 5527: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5528: 	jr	%ra
	-- is_outside.2834:
"10110000010111100000000000000000",	-- 5529: 	sf	%f2, [%sp + 0]
"10110000001111100000000000000001",	-- 5530: 	sf	%f1, [%sp + 1]
"00111100001111100000000000000010",	-- 5531: 	sw	%r1, [%sp + 2]
"10110000000111100000000000000011",	-- 5532: 	sf	%f0, [%sp + 3]
"00111111111111100000000000000100",	-- 5533: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5534: 	addi	%sp, %sp, 5
"01011000000000000000011001101001",	-- 5535: 	jal	o_param_x.2640
"10101011110111100000000000000101",	-- 5536: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5537: 	lw	%ra, [%sp + 4]
"10010011110000010000000000000011",	-- 5538: 	lf	%f1, [%sp + 3]
"11100100001000000000000000000000",	-- 5539: 	subf	%f0, %f1, %f0
"00111011110000010000000000000010",	-- 5540: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000100",	-- 5541: 	sf	%f0, [%sp + 4]
"00111111111111100000000000000101",	-- 5542: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5543: 	addi	%sp, %sp, 6
"01011000000000000000011001101110",	-- 5544: 	jal	o_param_y.2642
"10101011110111100000000000000110",	-- 5545: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5546: 	lw	%ra, [%sp + 5]
"10010011110000010000000000000001",	-- 5547: 	lf	%f1, [%sp + 1]
"11100100001000000000000000000000",	-- 5548: 	subf	%f0, %f1, %f0
"00111011110000010000000000000010",	-- 5549: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000101",	-- 5550: 	sf	%f0, [%sp + 5]
"00111111111111100000000000000110",	-- 5551: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5552: 	addi	%sp, %sp, 7
"01011000000000000000011001110011",	-- 5553: 	jal	o_param_z.2644
"10101011110111100000000000000111",	-- 5554: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5555: 	lw	%ra, [%sp + 6]
"10010011110000010000000000000000",	-- 5556: 	lf	%f1, [%sp + 0]
"11100100001000000000000000000000",	-- 5557: 	subf	%f0, %f1, %f0
"00111011110000010000000000000010",	-- 5558: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000110",	-- 5559: 	sf	%f0, [%sp + 6]
"00111111111111100000000000000111",	-- 5560: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 5561: 	addi	%sp, %sp, 8
"01011000000000000000011001010000",	-- 5562: 	jal	o_form.2624
"10101011110111100000000000001000",	-- 5563: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 5564: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000001",	-- 5565: 	lli	%r2, 1
"00101000001000100000000000000110",	-- 5566: 	bneq	%r1, %r2, bneq_else.9079
"10010011110000000000000000000100",	-- 5567: 	lf	%f0, [%sp + 4]
"10010011110000010000000000000101",	-- 5568: 	lf	%f1, [%sp + 5]
"10010011110000100000000000000110",	-- 5569: 	lf	%f2, [%sp + 6]
"00111011110000010000000000000010",	-- 5570: 	lw	%r1, [%sp + 2]
"01010100000000000001010011100111",	-- 5571: 	j	is_rect_outside.2819
	-- bneq_else.9079:
"11001100000000100000000000000010",	-- 5572: 	lli	%r2, 2
"00101000001000100000000000000110",	-- 5573: 	bneq	%r1, %r2, bneq_else.9080
"10010011110000000000000000000100",	-- 5574: 	lf	%f0, [%sp + 4]
"10010011110000010000000000000101",	-- 5575: 	lf	%f1, [%sp + 5]
"10010011110000100000000000000110",	-- 5576: 	lf	%f2, [%sp + 6]
"00111011110000010000000000000010",	-- 5577: 	lw	%r1, [%sp + 2]
"01010100000000000001010100111101",	-- 5578: 	j	is_plane_outside.2824
	-- bneq_else.9080:
"10010011110000000000000000000100",	-- 5579: 	lf	%f0, [%sp + 4]
"10010011110000010000000000000101",	-- 5580: 	lf	%f1, [%sp + 5]
"10010011110000100000000000000110",	-- 5581: 	lf	%f2, [%sp + 6]
"00111011110000010000000000000010",	-- 5582: 	lw	%r1, [%sp + 2]
"01010100000000000001010101101001",	-- 5583: 	j	is_second_outside.2829
	-- check_all_inside.2839:
"00111011011000110000000000000001",	-- 5584: 	lw	%r3, [%r27 + 1]
"10000100010000010010000000000000",	-- 5585: 	add	%r4, %r2, %r1
"00111000100001000000000000000000",	-- 5586: 	lw	%r4, [%r4 + 0]
"11001100000001011111111111111111",	-- 5587: 	lli	%r5, -1
"11001000000001011111111111111111",	-- 5588: 	lhi	%r5, -1
"00101000100001010000000000000011",	-- 5589: 	bneq	%r4, %r5, bneq_else.9081
"11001100000000010000000000000001",	-- 5590: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5591: 	jr	%ra
	-- bneq_else.9081:
"10000100011001000001100000000000",	-- 5592: 	add	%r3, %r3, %r4
"00111000011000110000000000000000",	-- 5593: 	lw	%r3, [%r3 + 0]
"10110000010111100000000000000000",	-- 5594: 	sf	%f2, [%sp + 0]
"10110000001111100000000000000001",	-- 5595: 	sf	%f1, [%sp + 1]
"10110000000111100000000000000010",	-- 5596: 	sf	%f0, [%sp + 2]
"00111100010111100000000000000011",	-- 5597: 	sw	%r2, [%sp + 3]
"00111111011111100000000000000100",	-- 5598: 	sw	%r27, [%sp + 4]
"00111100001111100000000000000101",	-- 5599: 	sw	%r1, [%sp + 5]
"10000100000000110000100000000000",	-- 5600: 	add	%r1, %r0, %r3
"00111111111111100000000000000110",	-- 5601: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5602: 	addi	%sp, %sp, 7
"01011000000000000001010110011001",	-- 5603: 	jal	is_outside.2834
"10101011110111100000000000000111",	-- 5604: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5605: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5606: 	lli	%r2, 0
"00101000001000100000000000001011",	-- 5607: 	bneq	%r1, %r2, bneq_else.9082
"11001100000000010000000000000001",	-- 5608: 	lli	%r1, 1
"00111011110000100000000000000101",	-- 5609: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 5610: 	add	%r1, %r2, %r1
"10010011110000000000000000000010",	-- 5611: 	lf	%f0, [%sp + 2]
"10010011110000010000000000000001",	-- 5612: 	lf	%f1, [%sp + 1]
"10010011110000100000000000000000",	-- 5613: 	lf	%f2, [%sp + 0]
"00111011110000100000000000000011",	-- 5614: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000100",	-- 5615: 	lw	%r27, [%sp + 4]
"00111011011110100000000000000000",	-- 5616: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5617: 	jr	%r26
	-- bneq_else.9082:
"11001100000000010000000000000000",	-- 5618: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5619: 	jr	%ra
	-- shadow_check_and_group.2845:
"00111011011000110000000000000111",	-- 5620: 	lw	%r3, [%r27 + 7]
"00111011011001000000000000000110",	-- 5621: 	lw	%r4, [%r27 + 6]
"00111011011001010000000000000101",	-- 5622: 	lw	%r5, [%r27 + 5]
"00111011011001100000000000000100",	-- 5623: 	lw	%r6, [%r27 + 4]
"00111011011001110000000000000011",	-- 5624: 	lw	%r7, [%r27 + 3]
"00111011011010000000000000000010",	-- 5625: 	lw	%r8, [%r27 + 2]
"00111011011010010000000000000001",	-- 5626: 	lw	%r9, [%r27 + 1]
"10000100010000010101000000000000",	-- 5627: 	add	%r10, %r2, %r1
"00111001010010100000000000000000",	-- 5628: 	lw	%r10, [%r10 + 0]
"11001100000010111111111111111111",	-- 5629: 	lli	%r11, -1
"11001000000010111111111111111111",	-- 5630: 	lhi	%r11, -1
"00101001010010110000000000000011",	-- 5631: 	bneq	%r10, %r11, bneq_else.9083
"11001100000000010000000000000000",	-- 5632: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5633: 	jr	%ra
	-- bneq_else.9083:
"10000100010000010101000000000000",	-- 5634: 	add	%r10, %r2, %r1
"00111001010010100000000000000000",	-- 5635: 	lw	%r10, [%r10 + 0]
"00111101001111100000000000000000",	-- 5636: 	sw	%r9, [%sp + 0]
"00111101000111100000000000000001",	-- 5637: 	sw	%r8, [%sp + 1]
"00111100111111100000000000000010",	-- 5638: 	sw	%r7, [%sp + 2]
"00111100010111100000000000000011",	-- 5639: 	sw	%r2, [%sp + 3]
"00111111011111100000000000000100",	-- 5640: 	sw	%r27, [%sp + 4]
"00111100001111100000000000000101",	-- 5641: 	sw	%r1, [%sp + 5]
"00111101010111100000000000000110",	-- 5642: 	sw	%r10, [%sp + 6]
"00111100101111100000000000000111",	-- 5643: 	sw	%r5, [%sp + 7]
"00111100100111100000000000001000",	-- 5644: 	sw	%r4, [%sp + 8]
"10000100000001100001000000000000",	-- 5645: 	add	%r2, %r0, %r6
"10000100000010100000100000000000",	-- 5646: 	add	%r1, %r0, %r10
"10000100000000111101100000000000",	-- 5647: 	add	%r27, %r0, %r3
"10000100000010000001100000000000",	-- 5648: 	add	%r3, %r0, %r8
"00111111111111100000000000001001",	-- 5649: 	sw	%ra, [%sp + 9]
"00111011011110100000000000000000",	-- 5650: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001010",	-- 5651: 	addi	%sp, %sp, 10
"01010011010000000000000000000000",	-- 5652: 	jalr	%r26
"10101011110111100000000000001010",	-- 5653: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 5654: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000000",	-- 5655: 	lli	%r2, 0
"00111011110000110000000000001000",	-- 5656: 	lw	%r3, [%sp + 8]
"10000100011000100001000000000000",	-- 5657: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 5658: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000000",	-- 5659: 	lli	%r2, 0
"10110000000111100000000000001001",	-- 5660: 	sf	%f0, [%sp + 9]
"00101000001000100000000000000011",	-- 5661: 	bneq	%r1, %r2, bneq_else.9084
"11001100000000010000000000000000",	-- 5662: 	lli	%r1, 0
"01010100000000000001011000100111",	-- 5663: 	j	bneq_cont.9085
	-- bneq_else.9084:
"00010100000000011100110011001101",	-- 5664: 	llif	%f1, -0.200000
"00010000000000011011111001001100",	-- 5665: 	lhif	%f1, -0.200000
"00111111111111100000000000001010",	-- 5666: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 5667: 	addi	%sp, %sp, 11
"01011000000000000000010011110001",	-- 5668: 	jal	fless.2532
"10101011110111100000000000001011",	-- 5669: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 5670: 	lw	%ra, [%sp + 10]
	-- bneq_cont.9085:
"11001100000000100000000000000000",	-- 5671: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 5672: 	bneq	%r1, %r2, bneq_else.9086
"00111011110000010000000000000110",	-- 5673: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000111",	-- 5674: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 5675: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 5676: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001010",	-- 5677: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 5678: 	addi	%sp, %sp, 11
"01011000000000000000011001010100",	-- 5679: 	jal	o_isinvert.2628
"10101011110111100000000000001011",	-- 5680: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 5681: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 5682: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5683: 	bneq	%r1, %r2, bneq_else.9087
"11001100000000010000000000000000",	-- 5684: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5685: 	jr	%ra
	-- bneq_else.9087:
"11001100000000010000000000000001",	-- 5686: 	lli	%r1, 1
"00111011110000100000000000000101",	-- 5687: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 5688: 	add	%r1, %r2, %r1
"00111011110000100000000000000011",	-- 5689: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000100",	-- 5690: 	lw	%r27, [%sp + 4]
"00111011011110100000000000000000",	-- 5691: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5692: 	jr	%r26
	-- bneq_else.9086:
"00010100000000001101011100001010",	-- 5693: 	llif	%f0, 0.010000
"00010000000000000011110000100011",	-- 5694: 	lhif	%f0, 0.010000
"10010011110000010000000000001001",	-- 5695: 	lf	%f1, [%sp + 9]
"11100000001000000000000000000000",	-- 5696: 	addf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 5697: 	lli	%r1, 0
"00111011110000100000000000000010",	-- 5698: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 5699: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 5700: 	lf	%f1, [%r1 + 0]
"11101000001000000000100000000000",	-- 5701: 	mulf	%f1, %f1, %f0
"11001100000000010000000000000000",	-- 5702: 	lli	%r1, 0
"00111011110000110000000000000001",	-- 5703: 	lw	%r3, [%sp + 1]
"10000100011000010000100000000000",	-- 5704: 	add	%r1, %r3, %r1
"10010000001000100000000000000000",	-- 5705: 	lf	%f2, [%r1 + 0]
"11100000001000100000100000000000",	-- 5706: 	addf	%f1, %f1, %f2
"11001100000000010000000000000001",	-- 5707: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 5708: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 5709: 	lf	%f2, [%r1 + 0]
"11101000010000000001000000000000",	-- 5710: 	mulf	%f2, %f2, %f0
"11001100000000010000000000000001",	-- 5711: 	lli	%r1, 1
"10000100011000010000100000000000",	-- 5712: 	add	%r1, %r3, %r1
"10010000001000110000000000000000",	-- 5713: 	lf	%f3, [%r1 + 0]
"11100000010000110001000000000000",	-- 5714: 	addf	%f2, %f2, %f3
"11001100000000010000000000000010",	-- 5715: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 5716: 	add	%r1, %r2, %r1
"10010000001000110000000000000000",	-- 5717: 	lf	%f3, [%r1 + 0]
"11101000011000000000000000000000",	-- 5718: 	mulf	%f0, %f3, %f0
"11001100000000010000000000000010",	-- 5719: 	lli	%r1, 2
"10000100011000010000100000000000",	-- 5720: 	add	%r1, %r3, %r1
"10010000001000110000000000000000",	-- 5721: 	lf	%f3, [%r1 + 0]
"11100000000000110000000000000000",	-- 5722: 	addf	%f0, %f0, %f3
"11001100000000010000000000000000",	-- 5723: 	lli	%r1, 0
"00111011110000100000000000000011",	-- 5724: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000000",	-- 5725: 	lw	%r27, [%sp + 0]
"00001100010111110000000000000000",	-- 5726: 	movf	%f31, %f2
"00001100000000100000000000000000",	-- 5727: 	movf	%f2, %f0
"00001100001000000000000000000000",	-- 5728: 	movf	%f0, %f1
"00001111111000010000000000000000",	-- 5729: 	movf	%f1, %f31
"00111111111111100000000000001010",	-- 5730: 	sw	%ra, [%sp + 10]
"00111011011110100000000000000000",	-- 5731: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001011",	-- 5732: 	addi	%sp, %sp, 11
"01010011010000000000000000000000",	-- 5733: 	jalr	%r26
"10101011110111100000000000001011",	-- 5734: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 5735: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 5736: 	lli	%r2, 0
"00101000001000100000000000001000",	-- 5737: 	bneq	%r1, %r2, bneq_else.9088
"11001100000000010000000000000001",	-- 5738: 	lli	%r1, 1
"00111011110000100000000000000101",	-- 5739: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 5740: 	add	%r1, %r2, %r1
"00111011110000100000000000000011",	-- 5741: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000100",	-- 5742: 	lw	%r27, [%sp + 4]
"00111011011110100000000000000000",	-- 5743: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5744: 	jr	%r26
	-- bneq_else.9088:
"11001100000000010000000000000001",	-- 5745: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5746: 	jr	%ra
	-- shadow_check_one_or_group.2848:
"00111011011000110000000000000010",	-- 5747: 	lw	%r3, [%r27 + 2]
"00111011011001000000000000000001",	-- 5748: 	lw	%r4, [%r27 + 1]
"10000100010000010010100000000000",	-- 5749: 	add	%r5, %r2, %r1
"00111000101001010000000000000000",	-- 5750: 	lw	%r5, [%r5 + 0]
"11001100000001101111111111111111",	-- 5751: 	lli	%r6, -1
"11001000000001101111111111111111",	-- 5752: 	lhi	%r6, -1
"00101000101001100000000000000011",	-- 5753: 	bneq	%r5, %r6, bneq_else.9089
"11001100000000010000000000000000",	-- 5754: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5755: 	jr	%ra
	-- bneq_else.9089:
"10000100100001010010000000000000",	-- 5756: 	add	%r4, %r4, %r5
"00111000100001000000000000000000",	-- 5757: 	lw	%r4, [%r4 + 0]
"11001100000001010000000000000000",	-- 5758: 	lli	%r5, 0
"00111100010111100000000000000000",	-- 5759: 	sw	%r2, [%sp + 0]
"00111111011111100000000000000001",	-- 5760: 	sw	%r27, [%sp + 1]
"00111100001111100000000000000010",	-- 5761: 	sw	%r1, [%sp + 2]
"10000100000001000001000000000000",	-- 5762: 	add	%r2, %r0, %r4
"10000100000001010000100000000000",	-- 5763: 	add	%r1, %r0, %r5
"10000100000000111101100000000000",	-- 5764: 	add	%r27, %r0, %r3
"00111111111111100000000000000011",	-- 5765: 	sw	%ra, [%sp + 3]
"00111011011110100000000000000000",	-- 5766: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000100",	-- 5767: 	addi	%sp, %sp, 4
"01010011010000000000000000000000",	-- 5768: 	jalr	%r26
"10101011110111100000000000000100",	-- 5769: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 5770: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000000",	-- 5771: 	lli	%r2, 0
"00101000001000100000000000001000",	-- 5772: 	bneq	%r1, %r2, bneq_else.9090
"11001100000000010000000000000001",	-- 5773: 	lli	%r1, 1
"00111011110000100000000000000010",	-- 5774: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 5775: 	add	%r1, %r2, %r1
"00111011110000100000000000000000",	-- 5776: 	lw	%r2, [%sp + 0]
"00111011110110110000000000000001",	-- 5777: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 5778: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5779: 	jr	%r26
	-- bneq_else.9090:
"11001100000000010000000000000001",	-- 5780: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5781: 	jr	%ra
	-- shadow_check_one_or_matrix.2851:
"00111011011000110000000000000101",	-- 5782: 	lw	%r3, [%r27 + 5]
"00111011011001000000000000000100",	-- 5783: 	lw	%r4, [%r27 + 4]
"00111011011001010000000000000011",	-- 5784: 	lw	%r5, [%r27 + 3]
"00111011011001100000000000000010",	-- 5785: 	lw	%r6, [%r27 + 2]
"00111011011001110000000000000001",	-- 5786: 	lw	%r7, [%r27 + 1]
"10000100010000010100000000000000",	-- 5787: 	add	%r8, %r2, %r1
"00111001000010000000000000000000",	-- 5788: 	lw	%r8, [%r8 + 0]
"11001100000010010000000000000000",	-- 5789: 	lli	%r9, 0
"10000101000010010100100000000000",	-- 5790: 	add	%r9, %r8, %r9
"00111001001010010000000000000000",	-- 5791: 	lw	%r9, [%r9 + 0]
"11001100000010101111111111111111",	-- 5792: 	lli	%r10, -1
"11001000000010101111111111111111",	-- 5793: 	lhi	%r10, -1
"00101001001010100000000000000011",	-- 5794: 	bneq	%r9, %r10, bneq_else.9091
"11001100000000010000000000000000",	-- 5795: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5796: 	jr	%ra
	-- bneq_else.9091:
"11001100000010100000000001100011",	-- 5797: 	lli	%r10, 99
"00111101000111100000000000000000",	-- 5798: 	sw	%r8, [%sp + 0]
"00111100101111100000000000000001",	-- 5799: 	sw	%r5, [%sp + 1]
"00111100010111100000000000000010",	-- 5800: 	sw	%r2, [%sp + 2]
"00111111011111100000000000000011",	-- 5801: 	sw	%r27, [%sp + 3]
"00111100001111100000000000000100",	-- 5802: 	sw	%r1, [%sp + 4]
"00101001001010100000000000000011",	-- 5803: 	bneq	%r9, %r10, bneq_else.9092
"11001100000000010000000000000001",	-- 5804: 	lli	%r1, 1
"01010100000000000001011011011010",	-- 5805: 	j	bneq_cont.9093
	-- bneq_else.9092:
"00111100100111100000000000000101",	-- 5806: 	sw	%r4, [%sp + 5]
"10000100000001100001000000000000",	-- 5807: 	add	%r2, %r0, %r6
"10000100000010010000100000000000",	-- 5808: 	add	%r1, %r0, %r9
"10000100000000111101100000000000",	-- 5809: 	add	%r27, %r0, %r3
"10000100000001110001100000000000",	-- 5810: 	add	%r3, %r0, %r7
"00111111111111100000000000000110",	-- 5811: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 5812: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 5813: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 5814: 	jalr	%r26
"10101011110111100000000000000111",	-- 5815: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5816: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5817: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5818: 	bneq	%r1, %r2, bneq_else.9094
"11001100000000010000000000000000",	-- 5819: 	lli	%r1, 0
"01010100000000000001011011011010",	-- 5820: 	j	bneq_cont.9095
	-- bneq_else.9094:
"11001100000000010000000000000000",	-- 5821: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 5822: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 5823: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 5824: 	lf	%f0, [%r1 + 0]
"00010100000000011100110011001101",	-- 5825: 	llif	%f1, -0.100000
"00010000000000011011110111001100",	-- 5826: 	lhif	%f1, -0.100000
"00111111111111100000000000000110",	-- 5827: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5828: 	addi	%sp, %sp, 7
"01011000000000000000010011110001",	-- 5829: 	jal	fless.2532
"10101011110111100000000000000111",	-- 5830: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5831: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5832: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5833: 	bneq	%r1, %r2, bneq_else.9096
"11001100000000010000000000000000",	-- 5834: 	lli	%r1, 0
"01010100000000000001011011011010",	-- 5835: 	j	bneq_cont.9097
	-- bneq_else.9096:
"11001100000000010000000000000001",	-- 5836: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 5837: 	lw	%r2, [%sp + 0]
"00111011110110110000000000000001",	-- 5838: 	lw	%r27, [%sp + 1]
"00111111111111100000000000000110",	-- 5839: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 5840: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 5841: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 5842: 	jalr	%r26
"10101011110111100000000000000111",	-- 5843: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5844: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5845: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5846: 	bneq	%r1, %r2, bneq_else.9098
"11001100000000010000000000000000",	-- 5847: 	lli	%r1, 0
"01010100000000000001011011011010",	-- 5848: 	j	bneq_cont.9099
	-- bneq_else.9098:
"11001100000000010000000000000001",	-- 5849: 	lli	%r1, 1
	-- bneq_cont.9099:
	-- bneq_cont.9097:
	-- bneq_cont.9095:
	-- bneq_cont.9093:
"11001100000000100000000000000000",	-- 5850: 	lli	%r2, 0
"00101000001000100000000000001000",	-- 5851: 	bneq	%r1, %r2, bneq_else.9100
"11001100000000010000000000000001",	-- 5852: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 5853: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5854: 	add	%r1, %r2, %r1
"00111011110000100000000000000010",	-- 5855: 	lw	%r2, [%sp + 2]
"00111011110110110000000000000011",	-- 5856: 	lw	%r27, [%sp + 3]
"00111011011110100000000000000000",	-- 5857: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5858: 	jr	%r26
	-- bneq_else.9100:
"11001100000000010000000000000001",	-- 5859: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 5860: 	lw	%r2, [%sp + 0]
"00111011110110110000000000000001",	-- 5861: 	lw	%r27, [%sp + 1]
"00111111111111100000000000000110",	-- 5862: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 5863: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 5864: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 5865: 	jalr	%r26
"10101011110111100000000000000111",	-- 5866: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5867: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5868: 	lli	%r2, 0
"00101000001000100000000000001000",	-- 5869: 	bneq	%r1, %r2, bneq_else.9101
"11001100000000010000000000000001",	-- 5870: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 5871: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5872: 	add	%r1, %r2, %r1
"00111011110000100000000000000010",	-- 5873: 	lw	%r2, [%sp + 2]
"00111011110110110000000000000011",	-- 5874: 	lw	%r27, [%sp + 3]
"00111011011110100000000000000000",	-- 5875: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5876: 	jr	%r26
	-- bneq_else.9101:
"11001100000000010000000000000001",	-- 5877: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5878: 	jr	%ra
	-- solve_each_element.2854:
"00111011011001000000000000001001",	-- 5879: 	lw	%r4, [%r27 + 9]
"00111011011001010000000000001000",	-- 5880: 	lw	%r5, [%r27 + 8]
"00111011011001100000000000000111",	-- 5881: 	lw	%r6, [%r27 + 7]
"00111011011001110000000000000110",	-- 5882: 	lw	%r7, [%r27 + 6]
"00111011011010000000000000000101",	-- 5883: 	lw	%r8, [%r27 + 5]
"00111011011010010000000000000100",	-- 5884: 	lw	%r9, [%r27 + 4]
"00111011011010100000000000000011",	-- 5885: 	lw	%r10, [%r27 + 3]
"00111011011010110000000000000010",	-- 5886: 	lw	%r11, [%r27 + 2]
"00111011011011000000000000000001",	-- 5887: 	lw	%r12, [%r27 + 1]
"10000100010000010110100000000000",	-- 5888: 	add	%r13, %r2, %r1
"00111001101011010000000000000000",	-- 5889: 	lw	%r13, [%r13 + 0]
"11001100000011101111111111111111",	-- 5890: 	lli	%r14, -1
"11001000000011101111111111111111",	-- 5891: 	lhi	%r14, -1
"00101001101011100000000000000010",	-- 5892: 	bneq	%r13, %r14, bneq_else.9102
"01001111111000000000000000000000",	-- 5893: 	jr	%ra
	-- bneq_else.9102:
"00111101001111100000000000000000",	-- 5894: 	sw	%r9, [%sp + 0]
"00111101011111100000000000000001",	-- 5895: 	sw	%r11, [%sp + 1]
"00111101010111100000000000000010",	-- 5896: 	sw	%r10, [%sp + 2]
"00111101100111100000000000000011",	-- 5897: 	sw	%r12, [%sp + 3]
"00111100101111100000000000000100",	-- 5898: 	sw	%r5, [%sp + 4]
"00111100100111100000000000000101",	-- 5899: 	sw	%r4, [%sp + 5]
"00111100110111100000000000000110",	-- 5900: 	sw	%r6, [%sp + 6]
"00111100011111100000000000000111",	-- 5901: 	sw	%r3, [%sp + 7]
"00111100010111100000000000001000",	-- 5902: 	sw	%r2, [%sp + 8]
"00111111011111100000000000001001",	-- 5903: 	sw	%r27, [%sp + 9]
"00111100001111100000000000001010",	-- 5904: 	sw	%r1, [%sp + 10]
"00111101101111100000000000001011",	-- 5905: 	sw	%r13, [%sp + 11]
"00111101000111100000000000001100",	-- 5906: 	sw	%r8, [%sp + 12]
"10000100000000110001000000000000",	-- 5907: 	add	%r2, %r0, %r3
"10000100000011010000100000000000",	-- 5908: 	add	%r1, %r0, %r13
"10000100000001111101100000000000",	-- 5909: 	add	%r27, %r0, %r7
"10000100000001010001100000000000",	-- 5910: 	add	%r3, %r0, %r5
"00111111111111100000000000001101",	-- 5911: 	sw	%ra, [%sp + 13]
"00111011011110100000000000000000",	-- 5912: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001110",	-- 5913: 	addi	%sp, %sp, 14
"01010011010000000000000000000000",	-- 5914: 	jalr	%r26
"10101011110111100000000000001110",	-- 5915: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 5916: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 5917: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 5918: 	bneq	%r1, %r2, bneq_else.9104
"00111011110000010000000000001011",	-- 5919: 	lw	%r1, [%sp + 11]
"00111011110000100000000000001100",	-- 5920: 	lw	%r2, [%sp + 12]
"10000100010000010000100000000000",	-- 5921: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 5922: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001101",	-- 5923: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 5924: 	addi	%sp, %sp, 14
"01011000000000000000011001010100",	-- 5925: 	jal	o_isinvert.2628
"10101011110111100000000000001110",	-- 5926: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 5927: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 5928: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 5929: 	bneq	%r1, %r2, bneq_else.9105
"01001111111000000000000000000000",	-- 5930: 	jr	%ra
	-- bneq_else.9105:
"11001100000000010000000000000001",	-- 5931: 	lli	%r1, 1
"00111011110000100000000000001010",	-- 5932: 	lw	%r2, [%sp + 10]
"10000100010000010000100000000000",	-- 5933: 	add	%r1, %r2, %r1
"00111011110000100000000000001000",	-- 5934: 	lw	%r2, [%sp + 8]
"00111011110000110000000000000111",	-- 5935: 	lw	%r3, [%sp + 7]
"00111011110110110000000000001001",	-- 5936: 	lw	%r27, [%sp + 9]
"00111011011110100000000000000000",	-- 5937: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5938: 	jr	%r26
	-- bneq_else.9104:
"11001100000000100000000000000000",	-- 5939: 	lli	%r2, 0
"00111011110000110000000000000110",	-- 5940: 	lw	%r3, [%sp + 6]
"10000100011000100001000000000000",	-- 5941: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 5942: 	lf	%f1, [%r2 + 0]
"00010100000000000000000000000000",	-- 5943: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 5944: 	lhif	%f0, 0.000000
"00111100001111100000000000001101",	-- 5945: 	sw	%r1, [%sp + 13]
"10110000001111100000000000001110",	-- 5946: 	sf	%f1, [%sp + 14]
"00111111111111100000000000001111",	-- 5947: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 5948: 	addi	%sp, %sp, 16
"01011000000000000000010011110001",	-- 5949: 	jal	fless.2532
"10101011110111100000000000010000",	-- 5950: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 5951: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 5952: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 5953: 	bneq	%r1, %r2, bneq_else.9107
"01010100000000000001011110011010",	-- 5954: 	j	bneq_cont.9108
	-- bneq_else.9107:
"11001100000000010000000000000000",	-- 5955: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 5956: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 5957: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 5958: 	lf	%f1, [%r1 + 0]
"10010011110000000000000000001110",	-- 5959: 	lf	%f0, [%sp + 14]
"00111111111111100000000000001111",	-- 5960: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 5961: 	addi	%sp, %sp, 16
"01011000000000000000010011110001",	-- 5962: 	jal	fless.2532
"10101011110111100000000000010000",	-- 5963: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 5964: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 5965: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 5966: 	bneq	%r1, %r2, bneq_else.9109
"01010100000000000001011110011010",	-- 5967: 	j	bneq_cont.9110
	-- bneq_else.9109:
"00010100000000001101011100001010",	-- 5968: 	llif	%f0, 0.010000
"00010000000000000011110000100011",	-- 5969: 	lhif	%f0, 0.010000
"10010011110000010000000000001110",	-- 5970: 	lf	%f1, [%sp + 14]
"11100000001000000000000000000000",	-- 5971: 	addf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 5972: 	lli	%r1, 0
"00111011110000100000000000000111",	-- 5973: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 5974: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 5975: 	lf	%f1, [%r1 + 0]
"11101000001000000000100000000000",	-- 5976: 	mulf	%f1, %f1, %f0
"11001100000000010000000000000000",	-- 5977: 	lli	%r1, 0
"00111011110000110000000000000100",	-- 5978: 	lw	%r3, [%sp + 4]
"10000100011000010000100000000000",	-- 5979: 	add	%r1, %r3, %r1
"10010000001000100000000000000000",	-- 5980: 	lf	%f2, [%r1 + 0]
"11100000001000100000100000000000",	-- 5981: 	addf	%f1, %f1, %f2
"11001100000000010000000000000001",	-- 5982: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 5983: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 5984: 	lf	%f2, [%r1 + 0]
"11101000010000000001000000000000",	-- 5985: 	mulf	%f2, %f2, %f0
"11001100000000010000000000000001",	-- 5986: 	lli	%r1, 1
"10000100011000010000100000000000",	-- 5987: 	add	%r1, %r3, %r1
"10010000001000110000000000000000",	-- 5988: 	lf	%f3, [%r1 + 0]
"11100000010000110001000000000000",	-- 5989: 	addf	%f2, %f2, %f3
"11001100000000010000000000000010",	-- 5990: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 5991: 	add	%r1, %r2, %r1
"10010000001000110000000000000000",	-- 5992: 	lf	%f3, [%r1 + 0]
"11101000011000000001100000000000",	-- 5993: 	mulf	%f3, %f3, %f0
"11001100000000010000000000000010",	-- 5994: 	lli	%r1, 2
"10000100011000010000100000000000",	-- 5995: 	add	%r1, %r3, %r1
"10010000001001000000000000000000",	-- 5996: 	lf	%f4, [%r1 + 0]
"11100000011001000001100000000000",	-- 5997: 	addf	%f3, %f3, %f4
"11001100000000010000000000000000",	-- 5998: 	lli	%r1, 0
"00111011110000110000000000001000",	-- 5999: 	lw	%r3, [%sp + 8]
"00111011110110110000000000000011",	-- 6000: 	lw	%r27, [%sp + 3]
"10110000011111100000000000001111",	-- 6001: 	sf	%f3, [%sp + 15]
"10110000010111100000000000010000",	-- 6002: 	sf	%f2, [%sp + 16]
"10110000001111100000000000010001",	-- 6003: 	sf	%f1, [%sp + 17]
"10110000000111100000000000010010",	-- 6004: 	sf	%f0, [%sp + 18]
"10000100000000110001000000000000",	-- 6005: 	add	%r2, %r0, %r3
"00001100001000000000000000000000",	-- 6006: 	movf	%f0, %f1
"00001100010000010000000000000000",	-- 6007: 	movf	%f1, %f2
"00001100011000100000000000000000",	-- 6008: 	movf	%f2, %f3
"00111111111111100000000000010011",	-- 6009: 	sw	%ra, [%sp + 19]
"00111011011110100000000000000000",	-- 6010: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010100",	-- 6011: 	addi	%sp, %sp, 20
"01010011010000000000000000000000",	-- 6012: 	jalr	%r26
"10101011110111100000000000010100",	-- 6013: 	subi	%sp, %sp, 20
"00111011110111110000000000010011",	-- 6014: 	lw	%ra, [%sp + 19]
"11001100000000100000000000000000",	-- 6015: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6016: 	bneq	%r1, %r2, bneq_else.9111
"01010100000000000001011110011010",	-- 6017: 	j	bneq_cont.9112
	-- bneq_else.9111:
"11001100000000010000000000000000",	-- 6018: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 6019: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 6020: 	add	%r1, %r2, %r1
"10010011110000000000000000010010",	-- 6021: 	lf	%f0, [%sp + 18]
"10110000000000010000000000000000",	-- 6022: 	sf	%f0, [%r1 + 0]
"10010011110000000000000000010001",	-- 6023: 	lf	%f0, [%sp + 17]
"10010011110000010000000000010000",	-- 6024: 	lf	%f1, [%sp + 16]
"10010011110000100000000000001111",	-- 6025: 	lf	%f2, [%sp + 15]
"00111011110000010000000000000010",	-- 6026: 	lw	%r1, [%sp + 2]
"00111111111111100000000000010011",	-- 6027: 	sw	%ra, [%sp + 19]
"10100111110111100000000000010100",	-- 6028: 	addi	%sp, %sp, 20
"01011000000000000000010100100100",	-- 6029: 	jal	vecset.2576
"10101011110111100000000000010100",	-- 6030: 	subi	%sp, %sp, 20
"00111011110111110000000000010011",	-- 6031: 	lw	%ra, [%sp + 19]
"11001100000000010000000000000000",	-- 6032: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 6033: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 6034: 	add	%r1, %r2, %r1
"00111011110000100000000000001011",	-- 6035: 	lw	%r2, [%sp + 11]
"00111100010000010000000000000000",	-- 6036: 	sw	%r2, [%r1 + 0]
"11001100000000010000000000000000",	-- 6037: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 6038: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6039: 	add	%r1, %r2, %r1
"00111011110000100000000000001101",	-- 6040: 	lw	%r2, [%sp + 13]
"00111100010000010000000000000000",	-- 6041: 	sw	%r2, [%r1 + 0]
	-- bneq_cont.9112:
	-- bneq_cont.9110:
	-- bneq_cont.9108:
"11001100000000010000000000000001",	-- 6042: 	lli	%r1, 1
"00111011110000100000000000001010",	-- 6043: 	lw	%r2, [%sp + 10]
"10000100010000010000100000000000",	-- 6044: 	add	%r1, %r2, %r1
"00111011110000100000000000001000",	-- 6045: 	lw	%r2, [%sp + 8]
"00111011110000110000000000000111",	-- 6046: 	lw	%r3, [%sp + 7]
"00111011110110110000000000001001",	-- 6047: 	lw	%r27, [%sp + 9]
"00111011011110100000000000000000",	-- 6048: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6049: 	jr	%r26
	-- solve_one_or_network.2858:
"00111011011001000000000000000010",	-- 6050: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 6051: 	lw	%r5, [%r27 + 1]
"10000100010000010011000000000000",	-- 6052: 	add	%r6, %r2, %r1
"00111000110001100000000000000000",	-- 6053: 	lw	%r6, [%r6 + 0]
"11001100000001111111111111111111",	-- 6054: 	lli	%r7, -1
"11001000000001111111111111111111",	-- 6055: 	lhi	%r7, -1
"00101000110001110000000000000010",	-- 6056: 	bneq	%r6, %r7, bneq_else.9113
"01001111111000000000000000000000",	-- 6057: 	jr	%ra
	-- bneq_else.9113:
"10000100101001100010100000000000",	-- 6058: 	add	%r5, %r5, %r6
"00111000101001010000000000000000",	-- 6059: 	lw	%r5, [%r5 + 0]
"11001100000001100000000000000000",	-- 6060: 	lli	%r6, 0
"00111100011111100000000000000000",	-- 6061: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 6062: 	sw	%r2, [%sp + 1]
"00111111011111100000000000000010",	-- 6063: 	sw	%r27, [%sp + 2]
"00111100001111100000000000000011",	-- 6064: 	sw	%r1, [%sp + 3]
"10000100000001010001000000000000",	-- 6065: 	add	%r2, %r0, %r5
"10000100000001100000100000000000",	-- 6066: 	add	%r1, %r0, %r6
"10000100000001001101100000000000",	-- 6067: 	add	%r27, %r0, %r4
"00111111111111100000000000000100",	-- 6068: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 6069: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 6070: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 6071: 	jalr	%r26
"10101011110111100000000000000101",	-- 6072: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6073: 	lw	%ra, [%sp + 4]
"11001100000000010000000000000001",	-- 6074: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 6075: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 6076: 	add	%r1, %r2, %r1
"00111011110000100000000000000001",	-- 6077: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 6078: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000010",	-- 6079: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 6080: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6081: 	jr	%r26
	-- trace_or_matrix.2862:
"00111011011001000000000000000101",	-- 6082: 	lw	%r4, [%r27 + 5]
"00111011011001010000000000000100",	-- 6083: 	lw	%r5, [%r27 + 4]
"00111011011001100000000000000011",	-- 6084: 	lw	%r6, [%r27 + 3]
"00111011011001110000000000000010",	-- 6085: 	lw	%r7, [%r27 + 2]
"00111011011010000000000000000001",	-- 6086: 	lw	%r8, [%r27 + 1]
"10000100010000010100100000000000",	-- 6087: 	add	%r9, %r2, %r1
"00111001001010010000000000000000",	-- 6088: 	lw	%r9, [%r9 + 0]
"11001100000010100000000000000000",	-- 6089: 	lli	%r10, 0
"10000101001010100101000000000000",	-- 6090: 	add	%r10, %r9, %r10
"00111001010010100000000000000000",	-- 6091: 	lw	%r10, [%r10 + 0]
"11001100000010111111111111111111",	-- 6092: 	lli	%r11, -1
"11001000000010111111111111111111",	-- 6093: 	lhi	%r11, -1
"00101001010010110000000000000010",	-- 6094: 	bneq	%r10, %r11, bneq_else.9115
"01001111111000000000000000000000",	-- 6095: 	jr	%ra
	-- bneq_else.9115:
"11001100000010110000000001100011",	-- 6096: 	lli	%r11, 99
"00111100011111100000000000000000",	-- 6097: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 6098: 	sw	%r2, [%sp + 1]
"00111111011111100000000000000010",	-- 6099: 	sw	%r27, [%sp + 2]
"00111100001111100000000000000011",	-- 6100: 	sw	%r1, [%sp + 3]
"00101001010010110000000000001100",	-- 6101: 	bneq	%r10, %r11, bneq_else.9117
"11001100000001000000000000000001",	-- 6102: 	lli	%r4, 1
"10000100000010010001000000000000",	-- 6103: 	add	%r2, %r0, %r9
"10000100000001000000100000000000",	-- 6104: 	add	%r1, %r0, %r4
"10000100000010001101100000000000",	-- 6105: 	add	%r27, %r0, %r8
"00111111111111100000000000000100",	-- 6106: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 6107: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 6108: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 6109: 	jalr	%r26
"10101011110111100000000000000101",	-- 6110: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6111: 	lw	%ra, [%sp + 4]
"01010100000000000001100000001100",	-- 6112: 	j	bneq_cont.9118
	-- bneq_else.9117:
"00111101001111100000000000000100",	-- 6113: 	sw	%r9, [%sp + 4]
"00111101000111100000000000000101",	-- 6114: 	sw	%r8, [%sp + 5]
"00111100100111100000000000000110",	-- 6115: 	sw	%r4, [%sp + 6]
"00111100110111100000000000000111",	-- 6116: 	sw	%r6, [%sp + 7]
"10000100000000110001000000000000",	-- 6117: 	add	%r2, %r0, %r3
"10000100000010100000100000000000",	-- 6118: 	add	%r1, %r0, %r10
"10000100000001111101100000000000",	-- 6119: 	add	%r27, %r0, %r7
"10000100000001010001100000000000",	-- 6120: 	add	%r3, %r0, %r5
"00111111111111100000000000001000",	-- 6121: 	sw	%ra, [%sp + 8]
"00111011011110100000000000000000",	-- 6122: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001001",	-- 6123: 	addi	%sp, %sp, 9
"01010011010000000000000000000000",	-- 6124: 	jalr	%r26
"10101011110111100000000000001001",	-- 6125: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6126: 	lw	%ra, [%sp + 8]
"11001100000000100000000000000000",	-- 6127: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6128: 	bneq	%r1, %r2, bneq_else.9119
"01010100000000000001100000001100",	-- 6129: 	j	bneq_cont.9120
	-- bneq_else.9119:
"11001100000000010000000000000000",	-- 6130: 	lli	%r1, 0
"00111011110000100000000000000111",	-- 6131: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 6132: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 6133: 	lf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 6134: 	lli	%r1, 0
"00111011110000100000000000000110",	-- 6135: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 6136: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6137: 	lf	%f1, [%r1 + 0]
"00111111111111100000000000001000",	-- 6138: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 6139: 	addi	%sp, %sp, 9
"01011000000000000000010011110001",	-- 6140: 	jal	fless.2532
"10101011110111100000000000001001",	-- 6141: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6142: 	lw	%ra, [%sp + 8]
"11001100000000100000000000000000",	-- 6143: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6144: 	bneq	%r1, %r2, bneq_else.9121
"01010100000000000001100000001100",	-- 6145: 	j	bneq_cont.9122
	-- bneq_else.9121:
"11001100000000010000000000000001",	-- 6146: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 6147: 	lw	%r2, [%sp + 4]
"00111011110000110000000000000000",	-- 6148: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000101",	-- 6149: 	lw	%r27, [%sp + 5]
"00111111111111100000000000001000",	-- 6150: 	sw	%ra, [%sp + 8]
"00111011011110100000000000000000",	-- 6151: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001001",	-- 6152: 	addi	%sp, %sp, 9
"01010011010000000000000000000000",	-- 6153: 	jalr	%r26
"10101011110111100000000000001001",	-- 6154: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6155: 	lw	%ra, [%sp + 8]
	-- bneq_cont.9122:
	-- bneq_cont.9120:
	-- bneq_cont.9118:
"11001100000000010000000000000001",	-- 6156: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 6157: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 6158: 	add	%r1, %r2, %r1
"00111011110000100000000000000001",	-- 6159: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 6160: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000010",	-- 6161: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 6162: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6163: 	jr	%r26
	-- judge_intersection.2866:
"00111011011000100000000000000011",	-- 6164: 	lw	%r2, [%r27 + 3]
"00111011011000110000000000000010",	-- 6165: 	lw	%r3, [%r27 + 2]
"00111011011001000000000000000001",	-- 6166: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 6167: 	lli	%r5, 0
"00010100000000000110101100101000",	-- 6168: 	llif	%f0, 1000000000.000000
"00010000000000000100111001101110",	-- 6169: 	lhif	%f0, 1000000000.000000
"10000100011001010010100000000000",	-- 6170: 	add	%r5, %r3, %r5
"10110000000001010000000000000000",	-- 6171: 	sf	%f0, [%r5 + 0]
"11001100000001010000000000000000",	-- 6172: 	lli	%r5, 0
"11001100000001100000000000000000",	-- 6173: 	lli	%r6, 0
"10000100100001100010000000000000",	-- 6174: 	add	%r4, %r4, %r6
"00111000100001000000000000000000",	-- 6175: 	lw	%r4, [%r4 + 0]
"00111100011111100000000000000000",	-- 6176: 	sw	%r3, [%sp + 0]
"10000100000000010001100000000000",	-- 6177: 	add	%r3, %r0, %r1
"10000100000000101101100000000000",	-- 6178: 	add	%r27, %r0, %r2
"10000100000001000001000000000000",	-- 6179: 	add	%r2, %r0, %r4
"10000100000001010000100000000000",	-- 6180: 	add	%r1, %r0, %r5
"00111111111111100000000000000001",	-- 6181: 	sw	%ra, [%sp + 1]
"00111011011110100000000000000000",	-- 6182: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000010",	-- 6183: 	addi	%sp, %sp, 2
"01010011010000000000000000000000",	-- 6184: 	jalr	%r26
"10101011110111100000000000000010",	-- 6185: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 6186: 	lw	%ra, [%sp + 1]
"11001100000000010000000000000000",	-- 6187: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 6188: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6189: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6190: 	lf	%f1, [%r1 + 0]
"00010100000000001100110011001101",	-- 6191: 	llif	%f0, -0.100000
"00010000000000001011110111001100",	-- 6192: 	lhif	%f0, -0.100000
"10110000001111100000000000000001",	-- 6193: 	sf	%f1, [%sp + 1]
"00111111111111100000000000000010",	-- 6194: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 6195: 	addi	%sp, %sp, 3
"01011000000000000000010011110001",	-- 6196: 	jal	fless.2532
"10101011110111100000000000000011",	-- 6197: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 6198: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000000",	-- 6199: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 6200: 	bneq	%r1, %r2, bneq_else.9123
"11001100000000010000000000000000",	-- 6201: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 6202: 	jr	%ra
	-- bneq_else.9123:
"00010100000000011011110000100000",	-- 6203: 	llif	%f1, 100000000.000000
"00010000000000010100110010111110",	-- 6204: 	lhif	%f1, 100000000.000000
"10010011110000000000000000000001",	-- 6205: 	lf	%f0, [%sp + 1]
"01010100000000000000010011110001",	-- 6206: 	j	fless.2532
	-- solve_each_element_fast.2868:
"00111011011001000000000000001001",	-- 6207: 	lw	%r4, [%r27 + 9]
"00111011011001010000000000001000",	-- 6208: 	lw	%r5, [%r27 + 8]
"00111011011001100000000000000111",	-- 6209: 	lw	%r6, [%r27 + 7]
"00111011011001110000000000000110",	-- 6210: 	lw	%r7, [%r27 + 6]
"00111011011010000000000000000101",	-- 6211: 	lw	%r8, [%r27 + 5]
"00111011011010010000000000000100",	-- 6212: 	lw	%r9, [%r27 + 4]
"00111011011010100000000000000011",	-- 6213: 	lw	%r10, [%r27 + 3]
"00111011011010110000000000000010",	-- 6214: 	lw	%r11, [%r27 + 2]
"00111011011011000000000000000001",	-- 6215: 	lw	%r12, [%r27 + 1]
"00111101001111100000000000000000",	-- 6216: 	sw	%r9, [%sp + 0]
"00111101011111100000000000000001",	-- 6217: 	sw	%r11, [%sp + 1]
"00111101010111100000000000000010",	-- 6218: 	sw	%r10, [%sp + 2]
"00111101100111100000000000000011",	-- 6219: 	sw	%r12, [%sp + 3]
"00111100101111100000000000000100",	-- 6220: 	sw	%r5, [%sp + 4]
"00111100100111100000000000000101",	-- 6221: 	sw	%r4, [%sp + 5]
"00111100111111100000000000000110",	-- 6222: 	sw	%r7, [%sp + 6]
"00111111011111100000000000000111",	-- 6223: 	sw	%r27, [%sp + 7]
"00111101000111100000000000001000",	-- 6224: 	sw	%r8, [%sp + 8]
"00111100011111100000000000001001",	-- 6225: 	sw	%r3, [%sp + 9]
"00111100110111100000000000001010",	-- 6226: 	sw	%r6, [%sp + 10]
"00111100001111100000000000001011",	-- 6227: 	sw	%r1, [%sp + 11]
"00111100010111100000000000001100",	-- 6228: 	sw	%r2, [%sp + 12]
"10000100000000110000100000000000",	-- 6229: 	add	%r1, %r0, %r3
"00111111111111100000000000001101",	-- 6230: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 6231: 	addi	%sp, %sp, 14
"01011000000000000000011010111010",	-- 6232: 	jal	d_vec.2683
"10101011110111100000000000001110",	-- 6233: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 6234: 	lw	%ra, [%sp + 13]
"00111011110000100000000000001011",	-- 6235: 	lw	%r2, [%sp + 11]
"00111011110000110000000000001100",	-- 6236: 	lw	%r3, [%sp + 12]
"10000100011000100010000000000000",	-- 6237: 	add	%r4, %r3, %r2
"00111000100001000000000000000000",	-- 6238: 	lw	%r4, [%r4 + 0]
"11001100000001011111111111111111",	-- 6239: 	lli	%r5, -1
"11001000000001011111111111111111",	-- 6240: 	lhi	%r5, -1
"00101000100001010000000000000010",	-- 6241: 	bneq	%r4, %r5, bneq_else.9124
"01001111111000000000000000000000",	-- 6242: 	jr	%ra
	-- bneq_else.9124:
"00111011110001010000000000001001",	-- 6243: 	lw	%r5, [%sp + 9]
"00111011110110110000000000001010",	-- 6244: 	lw	%r27, [%sp + 10]
"00111100001111100000000000001101",	-- 6245: 	sw	%r1, [%sp + 13]
"00111100100111100000000000001110",	-- 6246: 	sw	%r4, [%sp + 14]
"10000100000001010001000000000000",	-- 6247: 	add	%r2, %r0, %r5
"10000100000001000000100000000000",	-- 6248: 	add	%r1, %r0, %r4
"00111111111111100000000000001111",	-- 6249: 	sw	%ra, [%sp + 15]
"00111011011110100000000000000000",	-- 6250: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010000",	-- 6251: 	addi	%sp, %sp, 16
"01010011010000000000000000000000",	-- 6252: 	jalr	%r26
"10101011110111100000000000010000",	-- 6253: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 6254: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 6255: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 6256: 	bneq	%r1, %r2, bneq_else.9126
"00111011110000010000000000001110",	-- 6257: 	lw	%r1, [%sp + 14]
"00111011110000100000000000001000",	-- 6258: 	lw	%r2, [%sp + 8]
"10000100010000010000100000000000",	-- 6259: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 6260: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001111",	-- 6261: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 6262: 	addi	%sp, %sp, 16
"01011000000000000000011001010100",	-- 6263: 	jal	o_isinvert.2628
"10101011110111100000000000010000",	-- 6264: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 6265: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 6266: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6267: 	bneq	%r1, %r2, bneq_else.9127
"01001111111000000000000000000000",	-- 6268: 	jr	%ra
	-- bneq_else.9127:
"11001100000000010000000000000001",	-- 6269: 	lli	%r1, 1
"00111011110000100000000000001011",	-- 6270: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 6271: 	add	%r1, %r2, %r1
"00111011110000100000000000001100",	-- 6272: 	lw	%r2, [%sp + 12]
"00111011110000110000000000001001",	-- 6273: 	lw	%r3, [%sp + 9]
"00111011110110110000000000000111",	-- 6274: 	lw	%r27, [%sp + 7]
"00111011011110100000000000000000",	-- 6275: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6276: 	jr	%r26
	-- bneq_else.9126:
"11001100000000100000000000000000",	-- 6277: 	lli	%r2, 0
"00111011110000110000000000000110",	-- 6278: 	lw	%r3, [%sp + 6]
"10000100011000100001000000000000",	-- 6279: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 6280: 	lf	%f1, [%r2 + 0]
"00010100000000000000000000000000",	-- 6281: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 6282: 	lhif	%f0, 0.000000
"00111100001111100000000000001111",	-- 6283: 	sw	%r1, [%sp + 15]
"10110000001111100000000000010000",	-- 6284: 	sf	%f1, [%sp + 16]
"00111111111111100000000000010001",	-- 6285: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 6286: 	addi	%sp, %sp, 18
"01011000000000000000010011110001",	-- 6287: 	jal	fless.2532
"10101011110111100000000000010010",	-- 6288: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 6289: 	lw	%ra, [%sp + 17]
"11001100000000100000000000000000",	-- 6290: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6291: 	bneq	%r1, %r2, bneq_else.9129
"01010100000000000001100011101011",	-- 6292: 	j	bneq_cont.9130
	-- bneq_else.9129:
"11001100000000010000000000000000",	-- 6293: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 6294: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 6295: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6296: 	lf	%f1, [%r1 + 0]
"10010011110000000000000000010000",	-- 6297: 	lf	%f0, [%sp + 16]
"00111111111111100000000000010001",	-- 6298: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 6299: 	addi	%sp, %sp, 18
"01011000000000000000010011110001",	-- 6300: 	jal	fless.2532
"10101011110111100000000000010010",	-- 6301: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 6302: 	lw	%ra, [%sp + 17]
"11001100000000100000000000000000",	-- 6303: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6304: 	bneq	%r1, %r2, bneq_else.9131
"01010100000000000001100011101011",	-- 6305: 	j	bneq_cont.9132
	-- bneq_else.9131:
"00010100000000001101011100001010",	-- 6306: 	llif	%f0, 0.010000
"00010000000000000011110000100011",	-- 6307: 	lhif	%f0, 0.010000
"10010011110000010000000000010000",	-- 6308: 	lf	%f1, [%sp + 16]
"11100000001000000000000000000000",	-- 6309: 	addf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 6310: 	lli	%r1, 0
"00111011110000100000000000001101",	-- 6311: 	lw	%r2, [%sp + 13]
"10000100010000010000100000000000",	-- 6312: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6313: 	lf	%f1, [%r1 + 0]
"11101000001000000000100000000000",	-- 6314: 	mulf	%f1, %f1, %f0
"11001100000000010000000000000000",	-- 6315: 	lli	%r1, 0
"00111011110000110000000000000100",	-- 6316: 	lw	%r3, [%sp + 4]
"10000100011000010000100000000000",	-- 6317: 	add	%r1, %r3, %r1
"10010000001000100000000000000000",	-- 6318: 	lf	%f2, [%r1 + 0]
"11100000001000100000100000000000",	-- 6319: 	addf	%f1, %f1, %f2
"11001100000000010000000000000001",	-- 6320: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 6321: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 6322: 	lf	%f2, [%r1 + 0]
"11101000010000000001000000000000",	-- 6323: 	mulf	%f2, %f2, %f0
"11001100000000010000000000000001",	-- 6324: 	lli	%r1, 1
"10000100011000010000100000000000",	-- 6325: 	add	%r1, %r3, %r1
"10010000001000110000000000000000",	-- 6326: 	lf	%f3, [%r1 + 0]
"11100000010000110001000000000000",	-- 6327: 	addf	%f2, %f2, %f3
"11001100000000010000000000000010",	-- 6328: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 6329: 	add	%r1, %r2, %r1
"10010000001000110000000000000000",	-- 6330: 	lf	%f3, [%r1 + 0]
"11101000011000000001100000000000",	-- 6331: 	mulf	%f3, %f3, %f0
"11001100000000010000000000000010",	-- 6332: 	lli	%r1, 2
"10000100011000010000100000000000",	-- 6333: 	add	%r1, %r3, %r1
"10010000001001000000000000000000",	-- 6334: 	lf	%f4, [%r1 + 0]
"11100000011001000001100000000000",	-- 6335: 	addf	%f3, %f3, %f4
"11001100000000010000000000000000",	-- 6336: 	lli	%r1, 0
"00111011110000100000000000001100",	-- 6337: 	lw	%r2, [%sp + 12]
"00111011110110110000000000000011",	-- 6338: 	lw	%r27, [%sp + 3]
"10110000011111100000000000010001",	-- 6339: 	sf	%f3, [%sp + 17]
"10110000010111100000000000010010",	-- 6340: 	sf	%f2, [%sp + 18]
"10110000001111100000000000010011",	-- 6341: 	sf	%f1, [%sp + 19]
"10110000000111100000000000010100",	-- 6342: 	sf	%f0, [%sp + 20]
"00001100001000000000000000000000",	-- 6343: 	movf	%f0, %f1
"00001100010000010000000000000000",	-- 6344: 	movf	%f1, %f2
"00001100011000100000000000000000",	-- 6345: 	movf	%f2, %f3
"00111111111111100000000000010101",	-- 6346: 	sw	%ra, [%sp + 21]
"00111011011110100000000000000000",	-- 6347: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010110",	-- 6348: 	addi	%sp, %sp, 22
"01010011010000000000000000000000",	-- 6349: 	jalr	%r26
"10101011110111100000000000010110",	-- 6350: 	subi	%sp, %sp, 22
"00111011110111110000000000010101",	-- 6351: 	lw	%ra, [%sp + 21]
"11001100000000100000000000000000",	-- 6352: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6353: 	bneq	%r1, %r2, bneq_else.9133
"01010100000000000001100011101011",	-- 6354: 	j	bneq_cont.9134
	-- bneq_else.9133:
"11001100000000010000000000000000",	-- 6355: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 6356: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 6357: 	add	%r1, %r2, %r1
"10010011110000000000000000010100",	-- 6358: 	lf	%f0, [%sp + 20]
"10110000000000010000000000000000",	-- 6359: 	sf	%f0, [%r1 + 0]
"10010011110000000000000000010011",	-- 6360: 	lf	%f0, [%sp + 19]
"10010011110000010000000000010010",	-- 6361: 	lf	%f1, [%sp + 18]
"10010011110000100000000000010001",	-- 6362: 	lf	%f2, [%sp + 17]
"00111011110000010000000000000010",	-- 6363: 	lw	%r1, [%sp + 2]
"00111111111111100000000000010101",	-- 6364: 	sw	%ra, [%sp + 21]
"10100111110111100000000000010110",	-- 6365: 	addi	%sp, %sp, 22
"01011000000000000000010100100100",	-- 6366: 	jal	vecset.2576
"10101011110111100000000000010110",	-- 6367: 	subi	%sp, %sp, 22
"00111011110111110000000000010101",	-- 6368: 	lw	%ra, [%sp + 21]
"11001100000000010000000000000000",	-- 6369: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 6370: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 6371: 	add	%r1, %r2, %r1
"00111011110000100000000000001110",	-- 6372: 	lw	%r2, [%sp + 14]
"00111100010000010000000000000000",	-- 6373: 	sw	%r2, [%r1 + 0]
"11001100000000010000000000000000",	-- 6374: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 6375: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6376: 	add	%r1, %r2, %r1
"00111011110000100000000000001111",	-- 6377: 	lw	%r2, [%sp + 15]
"00111100010000010000000000000000",	-- 6378: 	sw	%r2, [%r1 + 0]
	-- bneq_cont.9134:
	-- bneq_cont.9132:
	-- bneq_cont.9130:
"11001100000000010000000000000001",	-- 6379: 	lli	%r1, 1
"00111011110000100000000000001011",	-- 6380: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 6381: 	add	%r1, %r2, %r1
"00111011110000100000000000001100",	-- 6382: 	lw	%r2, [%sp + 12]
"00111011110000110000000000001001",	-- 6383: 	lw	%r3, [%sp + 9]
"00111011110110110000000000000111",	-- 6384: 	lw	%r27, [%sp + 7]
"00111011011110100000000000000000",	-- 6385: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6386: 	jr	%r26
	-- solve_one_or_network_fast.2872:
"00111011011001000000000000000010",	-- 6387: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 6388: 	lw	%r5, [%r27 + 1]
"10000100010000010011000000000000",	-- 6389: 	add	%r6, %r2, %r1
"00111000110001100000000000000000",	-- 6390: 	lw	%r6, [%r6 + 0]
"11001100000001111111111111111111",	-- 6391: 	lli	%r7, -1
"11001000000001111111111111111111",	-- 6392: 	lhi	%r7, -1
"00101000110001110000000000000010",	-- 6393: 	bneq	%r6, %r7, bneq_else.9135
"01001111111000000000000000000000",	-- 6394: 	jr	%ra
	-- bneq_else.9135:
"10000100101001100010100000000000",	-- 6395: 	add	%r5, %r5, %r6
"00111000101001010000000000000000",	-- 6396: 	lw	%r5, [%r5 + 0]
"11001100000001100000000000000000",	-- 6397: 	lli	%r6, 0
"00111100011111100000000000000000",	-- 6398: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 6399: 	sw	%r2, [%sp + 1]
"00111111011111100000000000000010",	-- 6400: 	sw	%r27, [%sp + 2]
"00111100001111100000000000000011",	-- 6401: 	sw	%r1, [%sp + 3]
"10000100000001010001000000000000",	-- 6402: 	add	%r2, %r0, %r5
"10000100000001100000100000000000",	-- 6403: 	add	%r1, %r0, %r6
"10000100000001001101100000000000",	-- 6404: 	add	%r27, %r0, %r4
"00111111111111100000000000000100",	-- 6405: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 6406: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 6407: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 6408: 	jalr	%r26
"10101011110111100000000000000101",	-- 6409: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6410: 	lw	%ra, [%sp + 4]
"11001100000000010000000000000001",	-- 6411: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 6412: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 6413: 	add	%r1, %r2, %r1
"00111011110000100000000000000001",	-- 6414: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 6415: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000010",	-- 6416: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 6417: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6418: 	jr	%r26
	-- trace_or_matrix_fast.2876:
"00111011011001000000000000000100",	-- 6419: 	lw	%r4, [%r27 + 4]
"00111011011001010000000000000011",	-- 6420: 	lw	%r5, [%r27 + 3]
"00111011011001100000000000000010",	-- 6421: 	lw	%r6, [%r27 + 2]
"00111011011001110000000000000001",	-- 6422: 	lw	%r7, [%r27 + 1]
"10000100010000010100000000000000",	-- 6423: 	add	%r8, %r2, %r1
"00111001000010000000000000000000",	-- 6424: 	lw	%r8, [%r8 + 0]
"11001100000010010000000000000000",	-- 6425: 	lli	%r9, 0
"10000101000010010100100000000000",	-- 6426: 	add	%r9, %r8, %r9
"00111001001010010000000000000000",	-- 6427: 	lw	%r9, [%r9 + 0]
"11001100000010101111111111111111",	-- 6428: 	lli	%r10, -1
"11001000000010101111111111111111",	-- 6429: 	lhi	%r10, -1
"00101001001010100000000000000010",	-- 6430: 	bneq	%r9, %r10, bneq_else.9137
"01001111111000000000000000000000",	-- 6431: 	jr	%ra
	-- bneq_else.9137:
"11001100000010100000000001100011",	-- 6432: 	lli	%r10, 99
"00111100011111100000000000000000",	-- 6433: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 6434: 	sw	%r2, [%sp + 1]
"00111111011111100000000000000010",	-- 6435: 	sw	%r27, [%sp + 2]
"00111100001111100000000000000011",	-- 6436: 	sw	%r1, [%sp + 3]
"00101001001010100000000000001100",	-- 6437: 	bneq	%r9, %r10, bneq_else.9139
"11001100000001000000000000000001",	-- 6438: 	lli	%r4, 1
"10000100000010000001000000000000",	-- 6439: 	add	%r2, %r0, %r8
"10000100000001000000100000000000",	-- 6440: 	add	%r1, %r0, %r4
"10000100000001111101100000000000",	-- 6441: 	add	%r27, %r0, %r7
"00111111111111100000000000000100",	-- 6442: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 6443: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 6444: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 6445: 	jalr	%r26
"10101011110111100000000000000101",	-- 6446: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6447: 	lw	%ra, [%sp + 4]
"01010100000000000001100101011011",	-- 6448: 	j	bneq_cont.9140
	-- bneq_else.9139:
"00111101000111100000000000000100",	-- 6449: 	sw	%r8, [%sp + 4]
"00111100111111100000000000000101",	-- 6450: 	sw	%r7, [%sp + 5]
"00111100100111100000000000000110",	-- 6451: 	sw	%r4, [%sp + 6]
"00111100110111100000000000000111",	-- 6452: 	sw	%r6, [%sp + 7]
"10000100000000110001000000000000",	-- 6453: 	add	%r2, %r0, %r3
"10000100000010010000100000000000",	-- 6454: 	add	%r1, %r0, %r9
"10000100000001011101100000000000",	-- 6455: 	add	%r27, %r0, %r5
"00111111111111100000000000001000",	-- 6456: 	sw	%ra, [%sp + 8]
"00111011011110100000000000000000",	-- 6457: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001001",	-- 6458: 	addi	%sp, %sp, 9
"01010011010000000000000000000000",	-- 6459: 	jalr	%r26
"10101011110111100000000000001001",	-- 6460: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6461: 	lw	%ra, [%sp + 8]
"11001100000000100000000000000000",	-- 6462: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6463: 	bneq	%r1, %r2, bneq_else.9141
"01010100000000000001100101011011",	-- 6464: 	j	bneq_cont.9142
	-- bneq_else.9141:
"11001100000000010000000000000000",	-- 6465: 	lli	%r1, 0
"00111011110000100000000000000111",	-- 6466: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 6467: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 6468: 	lf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 6469: 	lli	%r1, 0
"00111011110000100000000000000110",	-- 6470: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 6471: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6472: 	lf	%f1, [%r1 + 0]
"00111111111111100000000000001000",	-- 6473: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 6474: 	addi	%sp, %sp, 9
"01011000000000000000010011110001",	-- 6475: 	jal	fless.2532
"10101011110111100000000000001001",	-- 6476: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6477: 	lw	%ra, [%sp + 8]
"11001100000000100000000000000000",	-- 6478: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6479: 	bneq	%r1, %r2, bneq_else.9143
"01010100000000000001100101011011",	-- 6480: 	j	bneq_cont.9144
	-- bneq_else.9143:
"11001100000000010000000000000001",	-- 6481: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 6482: 	lw	%r2, [%sp + 4]
"00111011110000110000000000000000",	-- 6483: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000101",	-- 6484: 	lw	%r27, [%sp + 5]
"00111111111111100000000000001000",	-- 6485: 	sw	%ra, [%sp + 8]
"00111011011110100000000000000000",	-- 6486: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001001",	-- 6487: 	addi	%sp, %sp, 9
"01010011010000000000000000000000",	-- 6488: 	jalr	%r26
"10101011110111100000000000001001",	-- 6489: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6490: 	lw	%ra, [%sp + 8]
	-- bneq_cont.9144:
	-- bneq_cont.9142:
	-- bneq_cont.9140:
"11001100000000010000000000000001",	-- 6491: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 6492: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 6493: 	add	%r1, %r2, %r1
"00111011110000100000000000000001",	-- 6494: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 6495: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000010",	-- 6496: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 6497: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6498: 	jr	%r26
	-- judge_intersection_fast.2880:
"00111011011000100000000000000011",	-- 6499: 	lw	%r2, [%r27 + 3]
"00111011011000110000000000000010",	-- 6500: 	lw	%r3, [%r27 + 2]
"00111011011001000000000000000001",	-- 6501: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 6502: 	lli	%r5, 0
"00010100000000000110101100101000",	-- 6503: 	llif	%f0, 1000000000.000000
"00010000000000000100111001101110",	-- 6504: 	lhif	%f0, 1000000000.000000
"10000100011001010010100000000000",	-- 6505: 	add	%r5, %r3, %r5
"10110000000001010000000000000000",	-- 6506: 	sf	%f0, [%r5 + 0]
"11001100000001010000000000000000",	-- 6507: 	lli	%r5, 0
"11001100000001100000000000000000",	-- 6508: 	lli	%r6, 0
"10000100100001100010000000000000",	-- 6509: 	add	%r4, %r4, %r6
"00111000100001000000000000000000",	-- 6510: 	lw	%r4, [%r4 + 0]
"00111100011111100000000000000000",	-- 6511: 	sw	%r3, [%sp + 0]
"10000100000000010001100000000000",	-- 6512: 	add	%r3, %r0, %r1
"10000100000000101101100000000000",	-- 6513: 	add	%r27, %r0, %r2
"10000100000001000001000000000000",	-- 6514: 	add	%r2, %r0, %r4
"10000100000001010000100000000000",	-- 6515: 	add	%r1, %r0, %r5
"00111111111111100000000000000001",	-- 6516: 	sw	%ra, [%sp + 1]
"00111011011110100000000000000000",	-- 6517: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000010",	-- 6518: 	addi	%sp, %sp, 2
"01010011010000000000000000000000",	-- 6519: 	jalr	%r26
"10101011110111100000000000000010",	-- 6520: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 6521: 	lw	%ra, [%sp + 1]
"11001100000000010000000000000000",	-- 6522: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 6523: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6524: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6525: 	lf	%f1, [%r1 + 0]
"00010100000000001100110011001101",	-- 6526: 	llif	%f0, -0.100000
"00010000000000001011110111001100",	-- 6527: 	lhif	%f0, -0.100000
"10110000001111100000000000000001",	-- 6528: 	sf	%f1, [%sp + 1]
"00111111111111100000000000000010",	-- 6529: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 6530: 	addi	%sp, %sp, 3
"01011000000000000000010011110001",	-- 6531: 	jal	fless.2532
"10101011110111100000000000000011",	-- 6532: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 6533: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000000",	-- 6534: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 6535: 	bneq	%r1, %r2, bneq_else.9145
"11001100000000010000000000000000",	-- 6536: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 6537: 	jr	%ra
	-- bneq_else.9145:
"00010100000000011011110000100000",	-- 6538: 	llif	%f1, 100000000.000000
"00010000000000010100110010111110",	-- 6539: 	lhif	%f1, 100000000.000000
"10010011110000000000000000000001",	-- 6540: 	lf	%f0, [%sp + 1]
"01010100000000000000010011110001",	-- 6541: 	j	fless.2532
	-- get_nvector_rect.2882:
"00111011011000100000000000000010",	-- 6542: 	lw	%r2, [%r27 + 2]
"00111011011000110000000000000001",	-- 6543: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 6544: 	lli	%r4, 0
"10000100011001000001100000000000",	-- 6545: 	add	%r3, %r3, %r4
"00111000011000110000000000000000",	-- 6546: 	lw	%r3, [%r3 + 0]
"00111100010111100000000000000000",	-- 6547: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 6548: 	sw	%r1, [%sp + 1]
"00111100011111100000000000000010",	-- 6549: 	sw	%r3, [%sp + 2]
"10000100000000100000100000000000",	-- 6550: 	add	%r1, %r0, %r2
"00111111111111100000000000000011",	-- 6551: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 6552: 	addi	%sp, %sp, 4
"01011000000000000000010100111000",	-- 6553: 	jal	vecbzero.2584
"10101011110111100000000000000100",	-- 6554: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 6555: 	lw	%ra, [%sp + 3]
"11001100000000010000000000000001",	-- 6556: 	lli	%r1, 1
"00111011110000100000000000000010",	-- 6557: 	lw	%r2, [%sp + 2]
"10001000010000010000100000000000",	-- 6558: 	sub	%r1, %r2, %r1
"11001100000000110000000000000001",	-- 6559: 	lli	%r3, 1
"10001000010000110001000000000000",	-- 6560: 	sub	%r2, %r2, %r3
"00111011110000110000000000000001",	-- 6561: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 6562: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 6563: 	lf	%f0, [%r2 + 0]
"00111100001111100000000000000011",	-- 6564: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 6565: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 6566: 	addi	%sp, %sp, 5
"01011000000000000000010100000000",	-- 6567: 	jal	sgn.2568
"10101011110111100000000000000101",	-- 6568: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6569: 	lw	%ra, [%sp + 4]
"00111111111111100000000000000100",	-- 6570: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 6571: 	addi	%sp, %sp, 5
"01011000000000000010101001001111",	-- 6572: 	jal	yj_fneg
"10101011110111100000000000000101",	-- 6573: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6574: 	lw	%ra, [%sp + 4]
"00111011110000010000000000000011",	-- 6575: 	lw	%r1, [%sp + 3]
"00111011110000100000000000000000",	-- 6576: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6577: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6578: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 6579: 	jr	%ra
	-- get_nvector_plane.2884:
"00111011011000100000000000000001",	-- 6580: 	lw	%r2, [%r27 + 1]
"11001100000000110000000000000000",	-- 6581: 	lli	%r3, 0
"00111100001111100000000000000000",	-- 6582: 	sw	%r1, [%sp + 0]
"00111100011111100000000000000001",	-- 6583: 	sw	%r3, [%sp + 1]
"00111100010111100000000000000010",	-- 6584: 	sw	%r2, [%sp + 2]
"00111111111111100000000000000011",	-- 6585: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 6586: 	addi	%sp, %sp, 4
"01011000000000000000011001011000",	-- 6587: 	jal	o_param_a.2632
"10101011110111100000000000000100",	-- 6588: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 6589: 	lw	%ra, [%sp + 3]
"00111111111111100000000000000011",	-- 6590: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 6591: 	addi	%sp, %sp, 4
"01011000000000000010101001001111",	-- 6592: 	jal	yj_fneg
"10101011110111100000000000000100",	-- 6593: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 6594: 	lw	%ra, [%sp + 3]
"00111011110000010000000000000001",	-- 6595: 	lw	%r1, [%sp + 1]
"00111011110000100000000000000010",	-- 6596: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 6597: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6598: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 6599: 	lli	%r1, 1
"00111011110000110000000000000000",	-- 6600: 	lw	%r3, [%sp + 0]
"00111100001111100000000000000011",	-- 6601: 	sw	%r1, [%sp + 3]
"10000100000000110000100000000000",	-- 6602: 	add	%r1, %r0, %r3
"00111111111111100000000000000100",	-- 6603: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 6604: 	addi	%sp, %sp, 5
"01011000000000000000011001011101",	-- 6605: 	jal	o_param_b.2634
"10101011110111100000000000000101",	-- 6606: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6607: 	lw	%ra, [%sp + 4]
"00111111111111100000000000000100",	-- 6608: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 6609: 	addi	%sp, %sp, 5
"01011000000000000010101001001111",	-- 6610: 	jal	yj_fneg
"10101011110111100000000000000101",	-- 6611: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6612: 	lw	%ra, [%sp + 4]
"00111011110000010000000000000011",	-- 6613: 	lw	%r1, [%sp + 3]
"00111011110000100000000000000010",	-- 6614: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 6615: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6616: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 6617: 	lli	%r1, 2
"00111011110000110000000000000000",	-- 6618: 	lw	%r3, [%sp + 0]
"00111100001111100000000000000100",	-- 6619: 	sw	%r1, [%sp + 4]
"10000100000000110000100000000000",	-- 6620: 	add	%r1, %r0, %r3
"00111111111111100000000000000101",	-- 6621: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 6622: 	addi	%sp, %sp, 6
"01011000000000000000011001100010",	-- 6623: 	jal	o_param_c.2636
"10101011110111100000000000000110",	-- 6624: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 6625: 	lw	%ra, [%sp + 5]
"00111111111111100000000000000101",	-- 6626: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 6627: 	addi	%sp, %sp, 6
"01011000000000000010101001001111",	-- 6628: 	jal	yj_fneg
"10101011110111100000000000000110",	-- 6629: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 6630: 	lw	%ra, [%sp + 5]
"00111011110000010000000000000100",	-- 6631: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000010",	-- 6632: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 6633: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6634: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 6635: 	jr	%ra
	-- get_nvector_second.2886:
"00111011011000100000000000000010",	-- 6636: 	lw	%r2, [%r27 + 2]
"00111011011000110000000000000001",	-- 6637: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 6638: 	lli	%r4, 0
"10000100011001000010000000000000",	-- 6639: 	add	%r4, %r3, %r4
"10010000100000000000000000000000",	-- 6640: 	lf	%f0, [%r4 + 0]
"00111100010111100000000000000000",	-- 6641: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 6642: 	sw	%r1, [%sp + 1]
"00111100011111100000000000000010",	-- 6643: 	sw	%r3, [%sp + 2]
"10110000000111100000000000000011",	-- 6644: 	sf	%f0, [%sp + 3]
"00111111111111100000000000000100",	-- 6645: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 6646: 	addi	%sp, %sp, 5
"01011000000000000000011001101001",	-- 6647: 	jal	o_param_x.2640
"10101011110111100000000000000101",	-- 6648: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6649: 	lw	%ra, [%sp + 4]
"10010011110000010000000000000011",	-- 6650: 	lf	%f1, [%sp + 3]
"11100100001000000000000000000000",	-- 6651: 	subf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 6652: 	lli	%r1, 1
"00111011110000100000000000000010",	-- 6653: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 6654: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6655: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000001",	-- 6656: 	lw	%r1, [%sp + 1]
"10110000000111100000000000000100",	-- 6657: 	sf	%f0, [%sp + 4]
"10110000001111100000000000000101",	-- 6658: 	sf	%f1, [%sp + 5]
"00111111111111100000000000000110",	-- 6659: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 6660: 	addi	%sp, %sp, 7
"01011000000000000000011001101110",	-- 6661: 	jal	o_param_y.2642
"10101011110111100000000000000111",	-- 6662: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 6663: 	lw	%ra, [%sp + 6]
"10010011110000010000000000000101",	-- 6664: 	lf	%f1, [%sp + 5]
"11100100001000000000000000000000",	-- 6665: 	subf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 6666: 	lli	%r1, 2
"00111011110000100000000000000010",	-- 6667: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 6668: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6669: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000001",	-- 6670: 	lw	%r1, [%sp + 1]
"10110000000111100000000000000110",	-- 6671: 	sf	%f0, [%sp + 6]
"10110000001111100000000000000111",	-- 6672: 	sf	%f1, [%sp + 7]
"00111111111111100000000000001000",	-- 6673: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 6674: 	addi	%sp, %sp, 9
"01011000000000000000011001110011",	-- 6675: 	jal	o_param_z.2644
"10101011110111100000000000001001",	-- 6676: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6677: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000111",	-- 6678: 	lf	%f1, [%sp + 7]
"11100100001000000000000000000000",	-- 6679: 	subf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6680: 	lw	%r1, [%sp + 1]
"10110000000111100000000000001000",	-- 6681: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 6682: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 6683: 	addi	%sp, %sp, 10
"01011000000000000000011001011000",	-- 6684: 	jal	o_param_a.2632
"10101011110111100000000000001010",	-- 6685: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 6686: 	lw	%ra, [%sp + 9]
"10010011110000010000000000000100",	-- 6687: 	lf	%f1, [%sp + 4]
"11101000001000000000000000000000",	-- 6688: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6689: 	lw	%r1, [%sp + 1]
"10110000000111100000000000001001",	-- 6690: 	sf	%f0, [%sp + 9]
"00111111111111100000000000001010",	-- 6691: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 6692: 	addi	%sp, %sp, 11
"01011000000000000000011001011101",	-- 6693: 	jal	o_param_b.2634
"10101011110111100000000000001011",	-- 6694: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 6695: 	lw	%ra, [%sp + 10]
"10010011110000010000000000000110",	-- 6696: 	lf	%f1, [%sp + 6]
"11101000001000000000000000000000",	-- 6697: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6698: 	lw	%r1, [%sp + 1]
"10110000000111100000000000001010",	-- 6699: 	sf	%f0, [%sp + 10]
"00111111111111100000000000001011",	-- 6700: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 6701: 	addi	%sp, %sp, 12
"01011000000000000000011001100010",	-- 6702: 	jal	o_param_c.2636
"10101011110111100000000000001100",	-- 6703: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 6704: 	lw	%ra, [%sp + 11]
"10010011110000010000000000001000",	-- 6705: 	lf	%f1, [%sp + 8]
"11101000001000000000000000000000",	-- 6706: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6707: 	lw	%r1, [%sp + 1]
"10110000000111100000000000001011",	-- 6708: 	sf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 6709: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 6710: 	addi	%sp, %sp, 13
"01011000000000000000011001010110",	-- 6711: 	jal	o_isrot.2630
"10101011110111100000000000001101",	-- 6712: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 6713: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000000",	-- 6714: 	lli	%r2, 0
"00101000001000100000000000001111",	-- 6715: 	bneq	%r1, %r2, bneq_else.9148
"11001100000000010000000000000000",	-- 6716: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 6717: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6718: 	add	%r1, %r2, %r1
"10010011110000000000000000001001",	-- 6719: 	lf	%f0, [%sp + 9]
"10110000000000010000000000000000",	-- 6720: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 6721: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 6722: 	add	%r1, %r2, %r1
"10010011110000000000000000001010",	-- 6723: 	lf	%f0, [%sp + 10]
"10110000000000010000000000000000",	-- 6724: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 6725: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 6726: 	add	%r1, %r2, %r1
"10010011110000000000000000001011",	-- 6727: 	lf	%f0, [%sp + 11]
"10110000000000010000000000000000",	-- 6728: 	sf	%f0, [%r1 + 0]
"01010100000000000001101010101101",	-- 6729: 	j	bneq_cont.9149
	-- bneq_else.9148:
"11001100000000010000000000000000",	-- 6730: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 6731: 	lw	%r2, [%sp + 1]
"00111100001111100000000000001100",	-- 6732: 	sw	%r1, [%sp + 12]
"10000100000000100000100000000000",	-- 6733: 	add	%r1, %r0, %r2
"00111111111111100000000000001101",	-- 6734: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 6735: 	addi	%sp, %sp, 14
"01011000000000000000011010011011",	-- 6736: 	jal	o_param_r3.2660
"10101011110111100000000000001110",	-- 6737: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 6738: 	lw	%ra, [%sp + 13]
"10010011110000010000000000000110",	-- 6739: 	lf	%f1, [%sp + 6]
"11101000001000000000000000000000",	-- 6740: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6741: 	lw	%r1, [%sp + 1]
"10110000000111100000000000001101",	-- 6742: 	sf	%f0, [%sp + 13]
"00111111111111100000000000001110",	-- 6743: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 6744: 	addi	%sp, %sp, 15
"01011000000000000000011010010110",	-- 6745: 	jal	o_param_r2.2658
"10101011110111100000000000001111",	-- 6746: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 6747: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001000",	-- 6748: 	lf	%f1, [%sp + 8]
"11101000001000000000000000000000",	-- 6749: 	mulf	%f0, %f1, %f0
"10010011110000100000000000001101",	-- 6750: 	lf	%f2, [%sp + 13]
"11100000010000000000000000000000",	-- 6751: 	addf	%f0, %f2, %f0
"00111111111111100000000000001110",	-- 6752: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 6753: 	addi	%sp, %sp, 15
"01011000000000000000010011101011",	-- 6754: 	jal	fhalf.2528
"10101011110111100000000000001111",	-- 6755: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 6756: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001001",	-- 6757: 	lf	%f1, [%sp + 9]
"11100000001000000000000000000000",	-- 6758: 	addf	%f0, %f1, %f0
"00111011110000010000000000001100",	-- 6759: 	lw	%r1, [%sp + 12]
"00111011110000100000000000000000",	-- 6760: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6761: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6762: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 6763: 	lli	%r1, 1
"00111011110000110000000000000001",	-- 6764: 	lw	%r3, [%sp + 1]
"00111100001111100000000000001110",	-- 6765: 	sw	%r1, [%sp + 14]
"10000100000000110000100000000000",	-- 6766: 	add	%r1, %r0, %r3
"00111111111111100000000000001111",	-- 6767: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 6768: 	addi	%sp, %sp, 16
"01011000000000000000011010011011",	-- 6769: 	jal	o_param_r3.2660
"10101011110111100000000000010000",	-- 6770: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 6771: 	lw	%ra, [%sp + 15]
"10010011110000010000000000000100",	-- 6772: 	lf	%f1, [%sp + 4]
"11101000001000000000000000000000",	-- 6773: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6774: 	lw	%r1, [%sp + 1]
"10110000000111100000000000001111",	-- 6775: 	sf	%f0, [%sp + 15]
"00111111111111100000000000010000",	-- 6776: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 6777: 	addi	%sp, %sp, 17
"01011000000000000000011010010001",	-- 6778: 	jal	o_param_r1.2656
"10101011110111100000000000010001",	-- 6779: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 6780: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001000",	-- 6781: 	lf	%f1, [%sp + 8]
"11101000001000000000000000000000",	-- 6782: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001111",	-- 6783: 	lf	%f1, [%sp + 15]
"11100000001000000000000000000000",	-- 6784: 	addf	%f0, %f1, %f0
"00111111111111100000000000010000",	-- 6785: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 6786: 	addi	%sp, %sp, 17
"01011000000000000000010011101011",	-- 6787: 	jal	fhalf.2528
"10101011110111100000000000010001",	-- 6788: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 6789: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001010",	-- 6790: 	lf	%f1, [%sp + 10]
"11100000001000000000000000000000",	-- 6791: 	addf	%f0, %f1, %f0
"00111011110000010000000000001110",	-- 6792: 	lw	%r1, [%sp + 14]
"00111011110000100000000000000000",	-- 6793: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6794: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6795: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 6796: 	lli	%r1, 2
"00111011110000110000000000000001",	-- 6797: 	lw	%r3, [%sp + 1]
"00111100001111100000000000010000",	-- 6798: 	sw	%r1, [%sp + 16]
"10000100000000110000100000000000",	-- 6799: 	add	%r1, %r0, %r3
"00111111111111100000000000010001",	-- 6800: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 6801: 	addi	%sp, %sp, 18
"01011000000000000000011010010110",	-- 6802: 	jal	o_param_r2.2658
"10101011110111100000000000010010",	-- 6803: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 6804: 	lw	%ra, [%sp + 17]
"10010011110000010000000000000100",	-- 6805: 	lf	%f1, [%sp + 4]
"11101000001000000000000000000000",	-- 6806: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6807: 	lw	%r1, [%sp + 1]
"10110000000111100000000000010001",	-- 6808: 	sf	%f0, [%sp + 17]
"00111111111111100000000000010010",	-- 6809: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 6810: 	addi	%sp, %sp, 19
"01011000000000000000011010010001",	-- 6811: 	jal	o_param_r1.2656
"10101011110111100000000000010011",	-- 6812: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 6813: 	lw	%ra, [%sp + 18]
"10010011110000010000000000000110",	-- 6814: 	lf	%f1, [%sp + 6]
"11101000001000000000000000000000",	-- 6815: 	mulf	%f0, %f1, %f0
"10010011110000010000000000010001",	-- 6816: 	lf	%f1, [%sp + 17]
"11100000001000000000000000000000",	-- 6817: 	addf	%f0, %f1, %f0
"00111111111111100000000000010010",	-- 6818: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 6819: 	addi	%sp, %sp, 19
"01011000000000000000010011101011",	-- 6820: 	jal	fhalf.2528
"10101011110111100000000000010011",	-- 6821: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 6822: 	lw	%ra, [%sp + 18]
"10010011110000010000000000001011",	-- 6823: 	lf	%f1, [%sp + 11]
"11100000001000000000000000000000",	-- 6824: 	addf	%f0, %f1, %f0
"00111011110000010000000000010000",	-- 6825: 	lw	%r1, [%sp + 16]
"00111011110000100000000000000000",	-- 6826: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6827: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6828: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9149:
"00111011110000010000000000000001",	-- 6829: 	lw	%r1, [%sp + 1]
"00111111111111100000000000010010",	-- 6830: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 6831: 	addi	%sp, %sp, 19
"01011000000000000000011001010100",	-- 6832: 	jal	o_isinvert.2628
"10101011110111100000000000010011",	-- 6833: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 6834: 	lw	%ra, [%sp + 18]
"10000100000000010001000000000000",	-- 6835: 	add	%r2, %r0, %r1
"00111011110000010000000000000000",	-- 6836: 	lw	%r1, [%sp + 0]
"01010100000000000000010101001110",	-- 6837: 	j	vecunit_sgn.2594
	-- get_nvector.2888:
"00111011011000110000000000000011",	-- 6838: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 6839: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 6840: 	lw	%r5, [%r27 + 1]
"00111100011111100000000000000000",	-- 6841: 	sw	%r3, [%sp + 0]
"00111100001111100000000000000001",	-- 6842: 	sw	%r1, [%sp + 1]
"00111100101111100000000000000010",	-- 6843: 	sw	%r5, [%sp + 2]
"00111100010111100000000000000011",	-- 6844: 	sw	%r2, [%sp + 3]
"00111100100111100000000000000100",	-- 6845: 	sw	%r4, [%sp + 4]
"00111111111111100000000000000101",	-- 6846: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 6847: 	addi	%sp, %sp, 6
"01011000000000000000011001010000",	-- 6848: 	jal	o_form.2624
"10101011110111100000000000000110",	-- 6849: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 6850: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000001",	-- 6851: 	lli	%r2, 1
"00101000001000100000000000000101",	-- 6852: 	bneq	%r1, %r2, bneq_else.9150
"00111011110000010000000000000011",	-- 6853: 	lw	%r1, [%sp + 3]
"00111011110110110000000000000100",	-- 6854: 	lw	%r27, [%sp + 4]
"00111011011110100000000000000000",	-- 6855: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6856: 	jr	%r26
	-- bneq_else.9150:
"11001100000000100000000000000010",	-- 6857: 	lli	%r2, 2
"00101000001000100000000000000101",	-- 6858: 	bneq	%r1, %r2, bneq_else.9151
"00111011110000010000000000000001",	-- 6859: 	lw	%r1, [%sp + 1]
"00111011110110110000000000000010",	-- 6860: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 6861: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6862: 	jr	%r26
	-- bneq_else.9151:
"00111011110000010000000000000001",	-- 6863: 	lw	%r1, [%sp + 1]
"00111011110110110000000000000000",	-- 6864: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 6865: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6866: 	jr	%r26
	-- utexture.2891:
"00111011011000110000000000000001",	-- 6867: 	lw	%r3, [%r27 + 1]
"00111100010111100000000000000000",	-- 6868: 	sw	%r2, [%sp + 0]
"00111100011111100000000000000001",	-- 6869: 	sw	%r3, [%sp + 1]
"00111100001111100000000000000010",	-- 6870: 	sw	%r1, [%sp + 2]
"00111111111111100000000000000011",	-- 6871: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 6872: 	addi	%sp, %sp, 4
"01011000000000000000011001001110",	-- 6873: 	jal	o_texturetype.2622
"10101011110111100000000000000100",	-- 6874: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 6875: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000000",	-- 6876: 	lli	%r2, 0
"00111011110000110000000000000010",	-- 6877: 	lw	%r3, [%sp + 2]
"00111100001111100000000000000011",	-- 6878: 	sw	%r1, [%sp + 3]
"00111100010111100000000000000100",	-- 6879: 	sw	%r2, [%sp + 4]
"10000100000000110000100000000000",	-- 6880: 	add	%r1, %r0, %r3
"00111111111111100000000000000101",	-- 6881: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 6882: 	addi	%sp, %sp, 6
"01011000000000000000011010000010",	-- 6883: 	jal	o_color_red.2650
"10101011110111100000000000000110",	-- 6884: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 6885: 	lw	%ra, [%sp + 5]
"00111011110000010000000000000100",	-- 6886: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000001",	-- 6887: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 6888: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6889: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 6890: 	lli	%r1, 1
"00111011110000110000000000000010",	-- 6891: 	lw	%r3, [%sp + 2]
"00111100001111100000000000000101",	-- 6892: 	sw	%r1, [%sp + 5]
"10000100000000110000100000000000",	-- 6893: 	add	%r1, %r0, %r3
"00111111111111100000000000000110",	-- 6894: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 6895: 	addi	%sp, %sp, 7
"01011000000000000000011010000111",	-- 6896: 	jal	o_color_green.2652
"10101011110111100000000000000111",	-- 6897: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 6898: 	lw	%ra, [%sp + 6]
"00111011110000010000000000000101",	-- 6899: 	lw	%r1, [%sp + 5]
"00111011110000100000000000000001",	-- 6900: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 6901: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6902: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 6903: 	lli	%r1, 2
"00111011110000110000000000000010",	-- 6904: 	lw	%r3, [%sp + 2]
"00111100001111100000000000000110",	-- 6905: 	sw	%r1, [%sp + 6]
"10000100000000110000100000000000",	-- 6906: 	add	%r1, %r0, %r3
"00111111111111100000000000000111",	-- 6907: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 6908: 	addi	%sp, %sp, 8
"01011000000000000000011010001100",	-- 6909: 	jal	o_color_blue.2654
"10101011110111100000000000001000",	-- 6910: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 6911: 	lw	%ra, [%sp + 7]
"00111011110000010000000000000110",	-- 6912: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000001",	-- 6913: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 6914: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6915: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 6916: 	lli	%r1, 1
"00111011110000110000000000000011",	-- 6917: 	lw	%r3, [%sp + 3]
"00101000011000010000000001100000",	-- 6918: 	bneq	%r3, %r1, bneq_else.9152
"11001100000000010000000000000000",	-- 6919: 	lli	%r1, 0
"00111011110000110000000000000000",	-- 6920: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 6921: 	add	%r1, %r3, %r1
"10010000001000000000000000000000",	-- 6922: 	lf	%f0, [%r1 + 0]
"00111011110000010000000000000010",	-- 6923: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000111",	-- 6924: 	sf	%f0, [%sp + 7]
"00111111111111100000000000001000",	-- 6925: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 6926: 	addi	%sp, %sp, 9
"01011000000000000000011001101001",	-- 6927: 	jal	o_param_x.2640
"10101011110111100000000000001001",	-- 6928: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6929: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000111",	-- 6930: 	lf	%f1, [%sp + 7]
"11100100001000000000000000000000",	-- 6931: 	subf	%f0, %f1, %f0
"00010100000000011100110011001101",	-- 6932: 	llif	%f1, 0.050000
"00010000000000010011110101001100",	-- 6933: 	lhif	%f1, 0.050000
"11101000000000010000100000000000",	-- 6934: 	mulf	%f1, %f0, %f1
"10110000000111100000000000001000",	-- 6935: 	sf	%f0, [%sp + 8]
"00001100001000000000000000000000",	-- 6936: 	movf	%f0, %f1
"00111111111111100000000000001001",	-- 6937: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 6938: 	addi	%sp, %sp, 10
"01011000000000000010101000110000",	-- 6939: 	jal	yj_floor
"10101011110111100000000000001010",	-- 6940: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 6941: 	lw	%ra, [%sp + 9]
"00010100000000010000000000000000",	-- 6942: 	llif	%f1, 20.000000
"00010000000000010100000110100000",	-- 6943: 	lhif	%f1, 20.000000
"11101000000000010000000000000000",	-- 6944: 	mulf	%f0, %f0, %f1
"10010011110000010000000000001000",	-- 6945: 	lf	%f1, [%sp + 8]
"11100100001000000000000000000000",	-- 6946: 	subf	%f0, %f1, %f0
"00010100000000010000000000000000",	-- 6947: 	llif	%f1, 10.000000
"00010000000000010100000100100000",	-- 6948: 	lhif	%f1, 10.000000
"00111111111111100000000000001001",	-- 6949: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 6950: 	addi	%sp, %sp, 10
"01011000000000000000010011110001",	-- 6951: 	jal	fless.2532
"10101011110111100000000000001010",	-- 6952: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 6953: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000010",	-- 6954: 	lli	%r2, 2
"00111011110000110000000000000000",	-- 6955: 	lw	%r3, [%sp + 0]
"10000100011000100001000000000000",	-- 6956: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 6957: 	lf	%f0, [%r2 + 0]
"00111011110000100000000000000010",	-- 6958: 	lw	%r2, [%sp + 2]
"00111100001111100000000000001001",	-- 6959: 	sw	%r1, [%sp + 9]
"10110000000111100000000000001010",	-- 6960: 	sf	%f0, [%sp + 10]
"10000100000000100000100000000000",	-- 6961: 	add	%r1, %r0, %r2
"00111111111111100000000000001011",	-- 6962: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 6963: 	addi	%sp, %sp, 12
"01011000000000000000011001110011",	-- 6964: 	jal	o_param_z.2644
"10101011110111100000000000001100",	-- 6965: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 6966: 	lw	%ra, [%sp + 11]
"10010011110000010000000000001010",	-- 6967: 	lf	%f1, [%sp + 10]
"11100100001000000000000000000000",	-- 6968: 	subf	%f0, %f1, %f0
"00010100000000011100110011001101",	-- 6969: 	llif	%f1, 0.050000
"00010000000000010011110101001100",	-- 6970: 	lhif	%f1, 0.050000
"11101000000000010000100000000000",	-- 6971: 	mulf	%f1, %f0, %f1
"10110000000111100000000000001011",	-- 6972: 	sf	%f0, [%sp + 11]
"00001100001000000000000000000000",	-- 6973: 	movf	%f0, %f1
"00111111111111100000000000001100",	-- 6974: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 6975: 	addi	%sp, %sp, 13
"01011000000000000010101000110000",	-- 6976: 	jal	yj_floor
"10101011110111100000000000001101",	-- 6977: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 6978: 	lw	%ra, [%sp + 12]
"00010100000000010000000000000000",	-- 6979: 	llif	%f1, 20.000000
"00010000000000010100000110100000",	-- 6980: 	lhif	%f1, 20.000000
"11101000000000010000000000000000",	-- 6981: 	mulf	%f0, %f0, %f1
"10010011110000010000000000001011",	-- 6982: 	lf	%f1, [%sp + 11]
"11100100001000000000000000000000",	-- 6983: 	subf	%f0, %f1, %f0
"00010100000000010000000000000000",	-- 6984: 	llif	%f1, 10.000000
"00010000000000010100000100100000",	-- 6985: 	lhif	%f1, 10.000000
"00111111111111100000000000001100",	-- 6986: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 6987: 	addi	%sp, %sp, 13
"01011000000000000000010011110001",	-- 6988: 	jal	fless.2532
"10101011110111100000000000001101",	-- 6989: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 6990: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000001",	-- 6991: 	lli	%r2, 1
"11001100000000110000000000000000",	-- 6992: 	lli	%r3, 0
"00111011110001000000000000001001",	-- 6993: 	lw	%r4, [%sp + 9]
"00101000100000110000000000001001",	-- 6994: 	bneq	%r4, %r3, bneq_else.9153
"11001100000000110000000000000000",	-- 6995: 	lli	%r3, 0
"00101000001000110000000000000100",	-- 6996: 	bneq	%r1, %r3, bneq_else.9155
"00010100000000000000000000000000",	-- 6997: 	llif	%f0, 255.000000
"00010000000000000100001101111111",	-- 6998: 	lhif	%f0, 255.000000
"01010100000000000001101101011010",	-- 6999: 	j	bneq_cont.9156
	-- bneq_else.9155:
"00010100000000000000000000000000",	-- 7000: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 7001: 	lhif	%f0, 0.000000
	-- bneq_cont.9156:
"01010100000000000001101101100010",	-- 7002: 	j	bneq_cont.9154
	-- bneq_else.9153:
"11001100000000110000000000000000",	-- 7003: 	lli	%r3, 0
"00101000001000110000000000000100",	-- 7004: 	bneq	%r1, %r3, bneq_else.9157
"00010100000000000000000000000000",	-- 7005: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 7006: 	lhif	%f0, 0.000000
"01010100000000000001101101100010",	-- 7007: 	j	bneq_cont.9158
	-- bneq_else.9157:
"00010100000000000000000000000000",	-- 7008: 	llif	%f0, 255.000000
"00010000000000000100001101111111",	-- 7009: 	lhif	%f0, 255.000000
	-- bneq_cont.9158:
	-- bneq_cont.9154:
"00111011110000010000000000000001",	-- 7010: 	lw	%r1, [%sp + 1]
"10000100001000100000100000000000",	-- 7011: 	add	%r1, %r1, %r2
"10110000000000010000000000000000",	-- 7012: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 7013: 	jr	%ra
	-- bneq_else.9152:
"11001100000000010000000000000010",	-- 7014: 	lli	%r1, 2
"00101000011000010000000000100011",	-- 7015: 	bneq	%r3, %r1, bneq_else.9160
"11001100000000010000000000000001",	-- 7016: 	lli	%r1, 1
"00111011110000110000000000000000",	-- 7017: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 7018: 	add	%r1, %r3, %r1
"10010000001000000000000000000000",	-- 7019: 	lf	%f0, [%r1 + 0]
"00010100000000010000000000000000",	-- 7020: 	llif	%f1, 0.250000
"00010000000000010011111010000000",	-- 7021: 	lhif	%f1, 0.250000
"11101000000000010000000000000000",	-- 7022: 	mulf	%f0, %f0, %f1
"00111111111111100000000000001100",	-- 7023: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 7024: 	addi	%sp, %sp, 13
"01011000000000000000010001010111",	-- 7025: 	jal	sin.2516
"10101011110111100000000000001101",	-- 7026: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 7027: 	lw	%ra, [%sp + 12]
"00111111111111100000000000001100",	-- 7028: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 7029: 	addi	%sp, %sp, 13
"01011000000000000000010011101111",	-- 7030: 	jal	fsqr.2530
"10101011110111100000000000001101",	-- 7031: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 7032: 	lw	%ra, [%sp + 12]
"11001100000000010000000000000000",	-- 7033: 	lli	%r1, 0
"00010100000000010000000000000000",	-- 7034: 	llif	%f1, 255.000000
"00010000000000010100001101111111",	-- 7035: 	lhif	%f1, 255.000000
"11101000001000000000100000000000",	-- 7036: 	mulf	%f1, %f1, %f0
"00111011110000100000000000000001",	-- 7037: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 7038: 	add	%r1, %r2, %r1
"10110000001000010000000000000000",	-- 7039: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000001",	-- 7040: 	lli	%r1, 1
"00010100000000010000000000000000",	-- 7041: 	llif	%f1, 255.000000
"00010000000000010100001101111111",	-- 7042: 	lhif	%f1, 255.000000
"00010100000000100000000000000000",	-- 7043: 	llif	%f2, 1.000000
"00010000000000100011111110000000",	-- 7044: 	lhif	%f2, 1.000000
"11100100010000000000000000000000",	-- 7045: 	subf	%f0, %f2, %f0
"11101000001000000000000000000000",	-- 7046: 	mulf	%f0, %f1, %f0
"10000100010000010000100000000000",	-- 7047: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 7048: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 7049: 	jr	%ra
	-- bneq_else.9160:
"11001100000000010000000000000011",	-- 7050: 	lli	%r1, 3
"00101000011000010000000001011100",	-- 7051: 	bneq	%r3, %r1, bneq_else.9162
"11001100000000010000000000000000",	-- 7052: 	lli	%r1, 0
"00111011110000110000000000000000",	-- 7053: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 7054: 	add	%r1, %r3, %r1
"10010000001000000000000000000000",	-- 7055: 	lf	%f0, [%r1 + 0]
"00111011110000010000000000000010",	-- 7056: 	lw	%r1, [%sp + 2]
"10110000000111100000000000001100",	-- 7057: 	sf	%f0, [%sp + 12]
"00111111111111100000000000001101",	-- 7058: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 7059: 	addi	%sp, %sp, 14
"01011000000000000000011001101001",	-- 7060: 	jal	o_param_x.2640
"10101011110111100000000000001110",	-- 7061: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 7062: 	lw	%ra, [%sp + 13]
"10010011110000010000000000001100",	-- 7063: 	lf	%f1, [%sp + 12]
"11100100001000000000000000000000",	-- 7064: 	subf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 7065: 	lli	%r1, 2
"00111011110000100000000000000000",	-- 7066: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 7067: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 7068: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000010",	-- 7069: 	lw	%r1, [%sp + 2]
"10110000000111100000000000001101",	-- 7070: 	sf	%f0, [%sp + 13]
"10110000001111100000000000001110",	-- 7071: 	sf	%f1, [%sp + 14]
"00111111111111100000000000001111",	-- 7072: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 7073: 	addi	%sp, %sp, 16
"01011000000000000000011001110011",	-- 7074: 	jal	o_param_z.2644
"10101011110111100000000000010000",	-- 7075: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 7076: 	lw	%ra, [%sp + 15]
"10010011110000010000000000001110",	-- 7077: 	lf	%f1, [%sp + 14]
"11100100001000000000000000000000",	-- 7078: 	subf	%f0, %f1, %f0
"10010011110000010000000000001101",	-- 7079: 	lf	%f1, [%sp + 13]
"10110000000111100000000000001111",	-- 7080: 	sf	%f0, [%sp + 15]
"00001100001000000000000000000000",	-- 7081: 	movf	%f0, %f1
"00111111111111100000000000010000",	-- 7082: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 7083: 	addi	%sp, %sp, 17
"01011000000000000000010011101111",	-- 7084: 	jal	fsqr.2530
"10101011110111100000000000010001",	-- 7085: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 7086: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001111",	-- 7087: 	lf	%f1, [%sp + 15]
"10110000000111100000000000010000",	-- 7088: 	sf	%f0, [%sp + 16]
"00001100001000000000000000000000",	-- 7089: 	movf	%f0, %f1
"00111111111111100000000000010001",	-- 7090: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 7091: 	addi	%sp, %sp, 18
"01011000000000000000010011101111",	-- 7092: 	jal	fsqr.2530
"10101011110111100000000000010010",	-- 7093: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 7094: 	lw	%ra, [%sp + 17]
"10010011110000010000000000010000",	-- 7095: 	lf	%f1, [%sp + 16]
"11100000001000000000000000000000",	-- 7096: 	addf	%f0, %f1, %f0
"00111111111111100000000000010001",	-- 7097: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 7098: 	addi	%sp, %sp, 18
"01011000000000000010101000101110",	-- 7099: 	jal	yj_sqrt
"10101011110111100000000000010010",	-- 7100: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 7101: 	lw	%ra, [%sp + 17]
"00010100000000010000000000000000",	-- 7102: 	llif	%f1, 10.000000
"00010000000000010100000100100000",	-- 7103: 	lhif	%f1, 10.000000
"11101100000000010000000000000000",	-- 7104: 	divf	%f0, %f0, %f1
"10110000000111100000000000010001",	-- 7105: 	sf	%f0, [%sp + 17]
"00111111111111100000000000010010",	-- 7106: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 7107: 	addi	%sp, %sp, 19
"01011000000000000010101000110000",	-- 7108: 	jal	yj_floor
"10101011110111100000000000010011",	-- 7109: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 7110: 	lw	%ra, [%sp + 18]
"10010011110000010000000000010001",	-- 7111: 	lf	%f1, [%sp + 17]
"11100100001000000000000000000000",	-- 7112: 	subf	%f0, %f1, %f0
"00010100000000010000111111011100",	-- 7113: 	llif	%f1, 3.141593
"00010000000000010100000001001001",	-- 7114: 	lhif	%f1, 3.141593
"11101000000000010000000000000000",	-- 7115: 	mulf	%f0, %f0, %f1
"00111111111111100000000000010010",	-- 7116: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 7117: 	addi	%sp, %sp, 19
"01011000000000000000010010010110",	-- 7118: 	jal	cos.2518
"10101011110111100000000000010011",	-- 7119: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 7120: 	lw	%ra, [%sp + 18]
"00111111111111100000000000010010",	-- 7121: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 7122: 	addi	%sp, %sp, 19
"01011000000000000000010011101111",	-- 7123: 	jal	fsqr.2530
"10101011110111100000000000010011",	-- 7124: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 7125: 	lw	%ra, [%sp + 18]
"11001100000000010000000000000001",	-- 7126: 	lli	%r1, 1
"00010100000000010000000000000000",	-- 7127: 	llif	%f1, 255.000000
"00010000000000010100001101111111",	-- 7128: 	lhif	%f1, 255.000000
"11101000000000010000100000000000",	-- 7129: 	mulf	%f1, %f0, %f1
"00111011110000100000000000000001",	-- 7130: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 7131: 	add	%r1, %r2, %r1
"10110000001000010000000000000000",	-- 7132: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 7133: 	lli	%r1, 2
"00010100000000010000000000000000",	-- 7134: 	llif	%f1, 1.000000
"00010000000000010011111110000000",	-- 7135: 	lhif	%f1, 1.000000
"11100100001000000000000000000000",	-- 7136: 	subf	%f0, %f1, %f0
"00010100000000010000000000000000",	-- 7137: 	llif	%f1, 255.000000
"00010000000000010100001101111111",	-- 7138: 	lhif	%f1, 255.000000
"11101000000000010000000000000000",	-- 7139: 	mulf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 7140: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 7141: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 7142: 	jr	%ra
	-- bneq_else.9162:
"11001100000000010000000000000100",	-- 7143: 	lli	%r1, 4
"00101000011000010000000011111000",	-- 7144: 	bneq	%r3, %r1, bneq_else.9164
"11001100000000010000000000000000",	-- 7145: 	lli	%r1, 0
"00111011110000110000000000000000",	-- 7146: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 7147: 	add	%r1, %r3, %r1
"10010000001000000000000000000000",	-- 7148: 	lf	%f0, [%r1 + 0]
"00111011110000010000000000000010",	-- 7149: 	lw	%r1, [%sp + 2]
"10110000000111100000000000010010",	-- 7150: 	sf	%f0, [%sp + 18]
"00111111111111100000000000010011",	-- 7151: 	sw	%ra, [%sp + 19]
"10100111110111100000000000010100",	-- 7152: 	addi	%sp, %sp, 20
"01011000000000000000011001101001",	-- 7153: 	jal	o_param_x.2640
"10101011110111100000000000010100",	-- 7154: 	subi	%sp, %sp, 20
"00111011110111110000000000010011",	-- 7155: 	lw	%ra, [%sp + 19]
"10010011110000010000000000010010",	-- 7156: 	lf	%f1, [%sp + 18]
"11100100001000000000000000000000",	-- 7157: 	subf	%f0, %f1, %f0
"00111011110000010000000000000010",	-- 7158: 	lw	%r1, [%sp + 2]
"10110000000111100000000000010011",	-- 7159: 	sf	%f0, [%sp + 19]
"00111111111111100000000000010100",	-- 7160: 	sw	%ra, [%sp + 20]
"10100111110111100000000000010101",	-- 7161: 	addi	%sp, %sp, 21
"01011000000000000000011001011000",	-- 7162: 	jal	o_param_a.2632
"10101011110111100000000000010101",	-- 7163: 	subi	%sp, %sp, 21
"00111011110111110000000000010100",	-- 7164: 	lw	%ra, [%sp + 20]
"00111111111111100000000000010100",	-- 7165: 	sw	%ra, [%sp + 20]
"10100111110111100000000000010101",	-- 7166: 	addi	%sp, %sp, 21
"01011000000000000010101000101110",	-- 7167: 	jal	yj_sqrt
"10101011110111100000000000010101",	-- 7168: 	subi	%sp, %sp, 21
"00111011110111110000000000010100",	-- 7169: 	lw	%ra, [%sp + 20]
"10010011110000010000000000010011",	-- 7170: 	lf	%f1, [%sp + 19]
"11101000001000000000000000000000",	-- 7171: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 7172: 	lli	%r1, 2
"00111011110000100000000000000000",	-- 7173: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 7174: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 7175: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000010",	-- 7176: 	lw	%r1, [%sp + 2]
"10110000000111100000000000010100",	-- 7177: 	sf	%f0, [%sp + 20]
"10110000001111100000000000010101",	-- 7178: 	sf	%f1, [%sp + 21]
"00111111111111100000000000010110",	-- 7179: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 7180: 	addi	%sp, %sp, 23
"01011000000000000000011001110011",	-- 7181: 	jal	o_param_z.2644
"10101011110111100000000000010111",	-- 7182: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 7183: 	lw	%ra, [%sp + 22]
"10010011110000010000000000010101",	-- 7184: 	lf	%f1, [%sp + 21]
"11100100001000000000000000000000",	-- 7185: 	subf	%f0, %f1, %f0
"00111011110000010000000000000010",	-- 7186: 	lw	%r1, [%sp + 2]
"10110000000111100000000000010110",	-- 7187: 	sf	%f0, [%sp + 22]
"00111111111111100000000000010111",	-- 7188: 	sw	%ra, [%sp + 23]
"10100111110111100000000000011000",	-- 7189: 	addi	%sp, %sp, 24
"01011000000000000000011001100010",	-- 7190: 	jal	o_param_c.2636
"10101011110111100000000000011000",	-- 7191: 	subi	%sp, %sp, 24
"00111011110111110000000000010111",	-- 7192: 	lw	%ra, [%sp + 23]
"00111111111111100000000000010111",	-- 7193: 	sw	%ra, [%sp + 23]
"10100111110111100000000000011000",	-- 7194: 	addi	%sp, %sp, 24
"01011000000000000010101000101110",	-- 7195: 	jal	yj_sqrt
"10101011110111100000000000011000",	-- 7196: 	subi	%sp, %sp, 24
"00111011110111110000000000010111",	-- 7197: 	lw	%ra, [%sp + 23]
"10010011110000010000000000010110",	-- 7198: 	lf	%f1, [%sp + 22]
"11101000001000000000000000000000",	-- 7199: 	mulf	%f0, %f1, %f0
"10010011110000010000000000010100",	-- 7200: 	lf	%f1, [%sp + 20]
"10110000000111100000000000010111",	-- 7201: 	sf	%f0, [%sp + 23]
"00001100001000000000000000000000",	-- 7202: 	movf	%f0, %f1
"00111111111111100000000000011000",	-- 7203: 	sw	%ra, [%sp + 24]
"10100111110111100000000000011001",	-- 7204: 	addi	%sp, %sp, 25
"01011000000000000000010011101111",	-- 7205: 	jal	fsqr.2530
"10101011110111100000000000011001",	-- 7206: 	subi	%sp, %sp, 25
"00111011110111110000000000011000",	-- 7207: 	lw	%ra, [%sp + 24]
"10010011110000010000000000010111",	-- 7208: 	lf	%f1, [%sp + 23]
"10110000000111100000000000011000",	-- 7209: 	sf	%f0, [%sp + 24]
"00001100001000000000000000000000",	-- 7210: 	movf	%f0, %f1
"00111111111111100000000000011001",	-- 7211: 	sw	%ra, [%sp + 25]
"10100111110111100000000000011010",	-- 7212: 	addi	%sp, %sp, 26
"01011000000000000000010011101111",	-- 7213: 	jal	fsqr.2530
"10101011110111100000000000011010",	-- 7214: 	subi	%sp, %sp, 26
"00111011110111110000000000011001",	-- 7215: 	lw	%ra, [%sp + 25]
"10010011110000010000000000011000",	-- 7216: 	lf	%f1, [%sp + 24]
"11100000001000000000000000000000",	-- 7217: 	addf	%f0, %f1, %f0
"10010011110000010000000000010100",	-- 7218: 	lf	%f1, [%sp + 20]
"10110000000111100000000000011001",	-- 7219: 	sf	%f0, [%sp + 25]
"00001100001000000000000000000000",	-- 7220: 	movf	%f0, %f1
"00111111111111100000000000011010",	-- 7221: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 7222: 	addi	%sp, %sp, 27
"01011000000000000010101001001101",	-- 7223: 	jal	yj_fabs
"10101011110111100000000000011011",	-- 7224: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 7225: 	lw	%ra, [%sp + 26]
"00010100000000011011011100010111",	-- 7226: 	llif	%f1, 0.000100
"00010000000000010011100011010001",	-- 7227: 	lhif	%f1, 0.000100
"00111111111111100000000000011010",	-- 7228: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 7229: 	addi	%sp, %sp, 27
"01011000000000000000010011110001",	-- 7230: 	jal	fless.2532
"10101011110111100000000000011011",	-- 7231: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 7232: 	lw	%ra, [%sp + 26]
"11001100000000100000000000000000",	-- 7233: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 7234: 	bneq	%r1, %r2, bneq_else.9165
"10010011110000000000000000010100",	-- 7235: 	lf	%f0, [%sp + 20]
"10010011110000010000000000010111",	-- 7236: 	lf	%f1, [%sp + 23]
"11101100001000000000000000000000",	-- 7237: 	divf	%f0, %f1, %f0
"00111111111111100000000000011010",	-- 7238: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 7239: 	addi	%sp, %sp, 27
"01011000000000000010101001001101",	-- 7240: 	jal	yj_fabs
"10101011110111100000000000011011",	-- 7241: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 7242: 	lw	%ra, [%sp + 26]
"00111111111111100000000000011010",	-- 7243: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 7244: 	addi	%sp, %sp, 27
"01011000000000000000010010011100",	-- 7245: 	jal	atan.2520
"10101011110111100000000000011011",	-- 7246: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 7247: 	lw	%ra, [%sp + 26]
"00010100000000010000000000000000",	-- 7248: 	llif	%f1, 30.000000
"00010000000000010100000111110000",	-- 7249: 	lhif	%f1, 30.000000
"11101000000000010000000000000000",	-- 7250: 	mulf	%f0, %f0, %f1
"00010100000000010000111111011100",	-- 7251: 	llif	%f1, 3.141593
"00010000000000010100000001001001",	-- 7252: 	lhif	%f1, 3.141593
"11101100000000010000000000000000",	-- 7253: 	divf	%f0, %f0, %f1
"01010100000000000001110001011001",	-- 7254: 	j	bneq_cont.9166
	-- bneq_else.9165:
"00010100000000000000000000000000",	-- 7255: 	llif	%f0, 15.000000
"00010000000000000100000101110000",	-- 7256: 	lhif	%f0, 15.000000
	-- bneq_cont.9166:
"10110000000111100000000000011010",	-- 7257: 	sf	%f0, [%sp + 26]
"00111111111111100000000000011011",	-- 7258: 	sw	%ra, [%sp + 27]
"10100111110111100000000000011100",	-- 7259: 	addi	%sp, %sp, 28
"01011000000000000010101000110000",	-- 7260: 	jal	yj_floor
"10101011110111100000000000011100",	-- 7261: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 7262: 	lw	%ra, [%sp + 27]
"10010011110000010000000000011010",	-- 7263: 	lf	%f1, [%sp + 26]
"11100100001000000000000000000000",	-- 7264: 	subf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 7265: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 7266: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 7267: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 7268: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000010",	-- 7269: 	lw	%r1, [%sp + 2]
"10110000000111100000000000011011",	-- 7270: 	sf	%f0, [%sp + 27]
"10110000001111100000000000011100",	-- 7271: 	sf	%f1, [%sp + 28]
"00111111111111100000000000011101",	-- 7272: 	sw	%ra, [%sp + 29]
"10100111110111100000000000011110",	-- 7273: 	addi	%sp, %sp, 30
"01011000000000000000011001101110",	-- 7274: 	jal	o_param_y.2642
"10101011110111100000000000011110",	-- 7275: 	subi	%sp, %sp, 30
"00111011110111110000000000011101",	-- 7276: 	lw	%ra, [%sp + 29]
"10010011110000010000000000011100",	-- 7277: 	lf	%f1, [%sp + 28]
"11100100001000000000000000000000",	-- 7278: 	subf	%f0, %f1, %f0
"00111011110000010000000000000010",	-- 7279: 	lw	%r1, [%sp + 2]
"10110000000111100000000000011101",	-- 7280: 	sf	%f0, [%sp + 29]
"00111111111111100000000000011110",	-- 7281: 	sw	%ra, [%sp + 30]
"10100111110111100000000000011111",	-- 7282: 	addi	%sp, %sp, 31
"01011000000000000000011001011101",	-- 7283: 	jal	o_param_b.2634
"10101011110111100000000000011111",	-- 7284: 	subi	%sp, %sp, 31
"00111011110111110000000000011110",	-- 7285: 	lw	%ra, [%sp + 30]
"00111111111111100000000000011110",	-- 7286: 	sw	%ra, [%sp + 30]
"10100111110111100000000000011111",	-- 7287: 	addi	%sp, %sp, 31
"01011000000000000010101000101110",	-- 7288: 	jal	yj_sqrt
"10101011110111100000000000011111",	-- 7289: 	subi	%sp, %sp, 31
"00111011110111110000000000011110",	-- 7290: 	lw	%ra, [%sp + 30]
"10010011110000010000000000011101",	-- 7291: 	lf	%f1, [%sp + 29]
"11101000001000000000000000000000",	-- 7292: 	mulf	%f0, %f1, %f0
"10010011110000010000000000011001",	-- 7293: 	lf	%f1, [%sp + 25]
"10110000000111100000000000011110",	-- 7294: 	sf	%f0, [%sp + 30]
"00001100001000000000000000000000",	-- 7295: 	movf	%f0, %f1
"00111111111111100000000000011111",	-- 7296: 	sw	%ra, [%sp + 31]
"10100111110111100000000000100000",	-- 7297: 	addi	%sp, %sp, 32
"01011000000000000010101001001101",	-- 7298: 	jal	yj_fabs
"10101011110111100000000000100000",	-- 7299: 	subi	%sp, %sp, 32
"00111011110111110000000000011111",	-- 7300: 	lw	%ra, [%sp + 31]
"00010100000000011011011100010111",	-- 7301: 	llif	%f1, 0.000100
"00010000000000010011100011010001",	-- 7302: 	lhif	%f1, 0.000100
"00111111111111100000000000011111",	-- 7303: 	sw	%ra, [%sp + 31]
"10100111110111100000000000100000",	-- 7304: 	addi	%sp, %sp, 32
"01011000000000000000010011110001",	-- 7305: 	jal	fless.2532
"10101011110111100000000000100000",	-- 7306: 	subi	%sp, %sp, 32
"00111011110111110000000000011111",	-- 7307: 	lw	%ra, [%sp + 31]
"11001100000000100000000000000000",	-- 7308: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 7309: 	bneq	%r1, %r2, bneq_else.9167
"10010011110000000000000000011001",	-- 7310: 	lf	%f0, [%sp + 25]
"10010011110000010000000000011110",	-- 7311: 	lf	%f1, [%sp + 30]
"11101100001000000000000000000000",	-- 7312: 	divf	%f0, %f1, %f0
"00111111111111100000000000011111",	-- 7313: 	sw	%ra, [%sp + 31]
"10100111110111100000000000100000",	-- 7314: 	addi	%sp, %sp, 32
"01011000000000000010101001001101",	-- 7315: 	jal	yj_fabs
"10101011110111100000000000100000",	-- 7316: 	subi	%sp, %sp, 32
"00111011110111110000000000011111",	-- 7317: 	lw	%ra, [%sp + 31]
"00111111111111100000000000011111",	-- 7318: 	sw	%ra, [%sp + 31]
"10100111110111100000000000100000",	-- 7319: 	addi	%sp, %sp, 32
"01011000000000000000010010011100",	-- 7320: 	jal	atan.2520
"10101011110111100000000000100000",	-- 7321: 	subi	%sp, %sp, 32
"00111011110111110000000000011111",	-- 7322: 	lw	%ra, [%sp + 31]
"00010100000000010000000000000000",	-- 7323: 	llif	%f1, 30.000000
"00010000000000010100000111110000",	-- 7324: 	lhif	%f1, 30.000000
"11101000000000010000000000000000",	-- 7325: 	mulf	%f0, %f0, %f1
"00010100000000010000111111011100",	-- 7326: 	llif	%f1, 3.141593
"00010000000000010100000001001001",	-- 7327: 	lhif	%f1, 3.141593
"11101100000000010000000000000000",	-- 7328: 	divf	%f0, %f0, %f1
"01010100000000000001110010100100",	-- 7329: 	j	bneq_cont.9168
	-- bneq_else.9167:
"00010100000000000000000000000000",	-- 7330: 	llif	%f0, 15.000000
"00010000000000000100000101110000",	-- 7331: 	lhif	%f0, 15.000000
	-- bneq_cont.9168:
"10110000000111100000000000011111",	-- 7332: 	sf	%f0, [%sp + 31]
"00111111111111100000000000100000",	-- 7333: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 7334: 	addi	%sp, %sp, 33
"01011000000000000010101000110000",	-- 7335: 	jal	yj_floor
"10101011110111100000000000100001",	-- 7336: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7337: 	lw	%ra, [%sp + 32]
"10010011110000010000000000011111",	-- 7338: 	lf	%f1, [%sp + 31]
"11100100001000000000000000000000",	-- 7339: 	subf	%f0, %f1, %f0
"00010100000000011001100110011010",	-- 7340: 	llif	%f1, 0.150000
"00010000000000010011111000011001",	-- 7341: 	lhif	%f1, 0.150000
"00010100000000100000000000000000",	-- 7342: 	llif	%f2, 0.500000
"00010000000000100011111100000000",	-- 7343: 	lhif	%f2, 0.500000
"10010011110000110000000000011011",	-- 7344: 	lf	%f3, [%sp + 27]
"11100100010000110001000000000000",	-- 7345: 	subf	%f2, %f2, %f3
"10110000000111100000000000100000",	-- 7346: 	sf	%f0, [%sp + 32]
"10110000001111100000000000100001",	-- 7347: 	sf	%f1, [%sp + 33]
"00001100010000000000000000000000",	-- 7348: 	movf	%f0, %f2
"00111111111111100000000000100010",	-- 7349: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 7350: 	addi	%sp, %sp, 35
"01011000000000000000010011101111",	-- 7351: 	jal	fsqr.2530
"10101011110111100000000000100011",	-- 7352: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 7353: 	lw	%ra, [%sp + 34]
"10010011110000010000000000100001",	-- 7354: 	lf	%f1, [%sp + 33]
"11100100001000000000000000000000",	-- 7355: 	subf	%f0, %f1, %f0
"00010100000000010000000000000000",	-- 7356: 	llif	%f1, 0.500000
"00010000000000010011111100000000",	-- 7357: 	lhif	%f1, 0.500000
"10010011110000100000000000100000",	-- 7358: 	lf	%f2, [%sp + 32]
"11100100001000100000100000000000",	-- 7359: 	subf	%f1, %f1, %f2
"10110000000111100000000000100010",	-- 7360: 	sf	%f0, [%sp + 34]
"00001100001000000000000000000000",	-- 7361: 	movf	%f0, %f1
"00111111111111100000000000100011",	-- 7362: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 7363: 	addi	%sp, %sp, 36
"01011000000000000000010011101111",	-- 7364: 	jal	fsqr.2530
"10101011110111100000000000100100",	-- 7365: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 7366: 	lw	%ra, [%sp + 35]
"10010011110000010000000000100010",	-- 7367: 	lf	%f1, [%sp + 34]
"11100100001000000000000000000000",	-- 7368: 	subf	%f0, %f1, %f0
"10110000000111100000000000100011",	-- 7369: 	sf	%f0, [%sp + 35]
"00111111111111100000000000100100",	-- 7370: 	sw	%ra, [%sp + 36]
"10100111110111100000000000100101",	-- 7371: 	addi	%sp, %sp, 37
"01011000000000000000010011011011",	-- 7372: 	jal	fisneg.2524
"10101011110111100000000000100101",	-- 7373: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 7374: 	lw	%ra, [%sp + 36]
"11001100000000100000000000000000",	-- 7375: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 7376: 	bneq	%r1, %r2, bneq_else.9169
"10010011110000000000000000100011",	-- 7377: 	lf	%f0, [%sp + 35]
"01010100000000000001110011010101",	-- 7378: 	j	bneq_cont.9170
	-- bneq_else.9169:
"00010100000000000000000000000000",	-- 7379: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 7380: 	lhif	%f0, 0.000000
	-- bneq_cont.9170:
"11001100000000010000000000000010",	-- 7381: 	lli	%r1, 2
"00010100000000010000000000000000",	-- 7382: 	llif	%f1, 255.000000
"00010000000000010100001101111111",	-- 7383: 	lhif	%f1, 255.000000
"11101000001000000000000000000000",	-- 7384: 	mulf	%f0, %f1, %f0
"00010100000000011001100110011010",	-- 7385: 	llif	%f1, 0.300000
"00010000000000010011111010011001",	-- 7386: 	lhif	%f1, 0.300000
"11101100000000010000000000000000",	-- 7387: 	divf	%f0, %f0, %f1
"00111011110000100000000000000001",	-- 7388: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 7389: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 7390: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 7391: 	jr	%ra
	-- bneq_else.9164:
"01001111111000000000000000000000",	-- 7392: 	jr	%ra
	-- add_light.2894:
"00111011011000010000000000000010",	-- 7393: 	lw	%r1, [%r27 + 2]
"00111011011000100000000000000001",	-- 7394: 	lw	%r2, [%r27 + 1]
"10110000010111100000000000000000",	-- 7395: 	sf	%f2, [%sp + 0]
"10110000001111100000000000000001",	-- 7396: 	sf	%f1, [%sp + 1]
"10110000000111100000000000000010",	-- 7397: 	sf	%f0, [%sp + 2]
"00111100001111100000000000000011",	-- 7398: 	sw	%r1, [%sp + 3]
"00111100010111100000000000000100",	-- 7399: 	sw	%r2, [%sp + 4]
"00111111111111100000000000000101",	-- 7400: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 7401: 	addi	%sp, %sp, 6
"01011000000000000000010011010100",	-- 7402: 	jal	fispos.2522
"10101011110111100000000000000110",	-- 7403: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 7404: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000000",	-- 7405: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 7406: 	bneq	%r1, %r2, bneq_else.9173
"01010100000000000001110011111000",	-- 7407: 	j	bneq_cont.9174
	-- bneq_else.9173:
"10010011110000000000000000000010",	-- 7408: 	lf	%f0, [%sp + 2]
"00111011110000010000000000000100",	-- 7409: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000011",	-- 7410: 	lw	%r2, [%sp + 3]
"00111111111111100000000000000101",	-- 7411: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 7412: 	addi	%sp, %sp, 6
"01011000000000000000010111001100",	-- 7413: 	jal	vecaccum.2605
"10101011110111100000000000000110",	-- 7414: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 7415: 	lw	%ra, [%sp + 5]
	-- bneq_cont.9174:
"10010011110000000000000000000001",	-- 7416: 	lf	%f0, [%sp + 1]
"00111111111111100000000000000101",	-- 7417: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 7418: 	addi	%sp, %sp, 6
"01011000000000000000010011010100",	-- 7419: 	jal	fispos.2522
"10101011110111100000000000000110",	-- 7420: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 7421: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000000",	-- 7422: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 7423: 	bneq	%r1, %r2, bneq_else.9175
"01001111111000000000000000000000",	-- 7424: 	jr	%ra
	-- bneq_else.9175:
"10010011110000000000000000000001",	-- 7425: 	lf	%f0, [%sp + 1]
"00111111111111100000000000000101",	-- 7426: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 7427: 	addi	%sp, %sp, 6
"01011000000000000000010011101111",	-- 7428: 	jal	fsqr.2530
"10101011110111100000000000000110",	-- 7429: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 7430: 	lw	%ra, [%sp + 5]
"00111111111111100000000000000101",	-- 7431: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 7432: 	addi	%sp, %sp, 6
"01011000000000000000010011101111",	-- 7433: 	jal	fsqr.2530
"10101011110111100000000000000110",	-- 7434: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 7435: 	lw	%ra, [%sp + 5]
"10010011110000010000000000000000",	-- 7436: 	lf	%f1, [%sp + 0]
"11101000000000010000000000000000",	-- 7437: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000000",	-- 7438: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 7439: 	lli	%r2, 0
"00111011110000110000000000000100",	-- 7440: 	lw	%r3, [%sp + 4]
"10000100011000100001000000000000",	-- 7441: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 7442: 	lf	%f1, [%r2 + 0]
"11100000001000000000100000000000",	-- 7443: 	addf	%f1, %f1, %f0
"10000100011000010000100000000000",	-- 7444: 	add	%r1, %r3, %r1
"10110000001000010000000000000000",	-- 7445: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000001",	-- 7446: 	lli	%r1, 1
"11001100000000100000000000000001",	-- 7447: 	lli	%r2, 1
"10000100011000100001000000000000",	-- 7448: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 7449: 	lf	%f1, [%r2 + 0]
"11100000001000000000100000000000",	-- 7450: 	addf	%f1, %f1, %f0
"10000100011000010000100000000000",	-- 7451: 	add	%r1, %r3, %r1
"10110000001000010000000000000000",	-- 7452: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 7453: 	lli	%r1, 2
"11001100000000100000000000000010",	-- 7454: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 7455: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 7456: 	lf	%f1, [%r2 + 0]
"11100000001000000000000000000000",	-- 7457: 	addf	%f0, %f1, %f0
"10000100011000010000100000000000",	-- 7458: 	add	%r1, %r3, %r1
"10110000000000010000000000000000",	-- 7459: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 7460: 	jr	%ra
	-- trace_reflections.2898:
"00111011011000110000000000001000",	-- 7461: 	lw	%r3, [%r27 + 8]
"00111011011001000000000000000111",	-- 7462: 	lw	%r4, [%r27 + 7]
"00111011011001010000000000000110",	-- 7463: 	lw	%r5, [%r27 + 6]
"00111011011001100000000000000101",	-- 7464: 	lw	%r6, [%r27 + 5]
"00111011011001110000000000000100",	-- 7465: 	lw	%r7, [%r27 + 4]
"00111011011010000000000000000011",	-- 7466: 	lw	%r8, [%r27 + 3]
"00111011011010010000000000000010",	-- 7467: 	lw	%r9, [%r27 + 2]
"00111011011010100000000000000001",	-- 7468: 	lw	%r10, [%r27 + 1]
"11001100000010110000000000000000",	-- 7469: 	lli	%r11, 0
"00110001011000010000000010000001",	-- 7470: 	bgt	%r11, %r1, bgt_else.9178
"10000100100000010010000000000000",	-- 7471: 	add	%r4, %r4, %r1
"00111000100001000000000000000000",	-- 7472: 	lw	%r4, [%r4 + 0]
"00111111011111100000000000000000",	-- 7473: 	sw	%r27, [%sp + 0]
"00111100001111100000000000000001",	-- 7474: 	sw	%r1, [%sp + 1]
"10110000001111100000000000000010",	-- 7475: 	sf	%f1, [%sp + 2]
"00111101010111100000000000000011",	-- 7476: 	sw	%r10, [%sp + 3]
"00111100010111100000000000000100",	-- 7477: 	sw	%r2, [%sp + 4]
"10110000000111100000000000000101",	-- 7478: 	sf	%f0, [%sp + 5]
"00111100110111100000000000000110",	-- 7479: 	sw	%r6, [%sp + 6]
"00111100011111100000000000000111",	-- 7480: 	sw	%r3, [%sp + 7]
"00111100101111100000000000001000",	-- 7481: 	sw	%r5, [%sp + 8]
"00111100100111100000000000001001",	-- 7482: 	sw	%r4, [%sp + 9]
"00111101000111100000000000001010",	-- 7483: 	sw	%r8, [%sp + 10]
"00111101001111100000000000001011",	-- 7484: 	sw	%r9, [%sp + 11]
"00111100111111100000000000001100",	-- 7485: 	sw	%r7, [%sp + 12]
"10000100000001000000100000000000",	-- 7486: 	add	%r1, %r0, %r4
"00111111111111100000000000001101",	-- 7487: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 7488: 	addi	%sp, %sp, 14
"01011000000000000000011011000000",	-- 7489: 	jal	r_dvec.2689
"10101011110111100000000000001110",	-- 7490: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 7491: 	lw	%ra, [%sp + 13]
"00111011110110110000000000001100",	-- 7492: 	lw	%r27, [%sp + 12]
"00111100001111100000000000001101",	-- 7493: 	sw	%r1, [%sp + 13]
"00111111111111100000000000001110",	-- 7494: 	sw	%ra, [%sp + 14]
"00111011011110100000000000000000",	-- 7495: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001111",	-- 7496: 	addi	%sp, %sp, 15
"01010011010000000000000000000000",	-- 7497: 	jalr	%r26
"10101011110111100000000000001111",	-- 7498: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 7499: 	lw	%ra, [%sp + 14]
"11001100000000100000000000000000",	-- 7500: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 7501: 	bneq	%r1, %r2, bneq_else.9179
"01010100000000000001110110100110",	-- 7502: 	j	bneq_cont.9180
	-- bneq_else.9179:
"11001100000000010000000000000000",	-- 7503: 	lli	%r1, 0
"00111011110000100000000000001011",	-- 7504: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 7505: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 7506: 	lw	%r1, [%r1 + 0]
"11001100000000100000000000000100",	-- 7507: 	lli	%r2, 4
"10001100001000100000100000000000",	-- 7508: 	mul	%r1, %r1, %r2
"11001100000000100000000000000000",	-- 7509: 	lli	%r2, 0
"00111011110000110000000000001010",	-- 7510: 	lw	%r3, [%sp + 10]
"10000100011000100001000000000000",	-- 7511: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 7512: 	lw	%r2, [%r2 + 0]
"10000100001000100000100000000000",	-- 7513: 	add	%r1, %r1, %r2
"00111011110000100000000000001001",	-- 7514: 	lw	%r2, [%sp + 9]
"00111100001111100000000000001110",	-- 7515: 	sw	%r1, [%sp + 14]
"10000100000000100000100000000000",	-- 7516: 	add	%r1, %r0, %r2
"00111111111111100000000000001111",	-- 7517: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 7518: 	addi	%sp, %sp, 16
"01011000000000000000011010111110",	-- 7519: 	jal	r_surface_id.2687
"10101011110111100000000000010000",	-- 7520: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 7521: 	lw	%ra, [%sp + 15]
"00111011110000100000000000001110",	-- 7522: 	lw	%r2, [%sp + 14]
"00101000010000010000000001000011",	-- 7523: 	bneq	%r2, %r1, bneq_else.9181
"11001100000000010000000000000000",	-- 7524: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 7525: 	lli	%r2, 0
"00111011110000110000000000001000",	-- 7526: 	lw	%r3, [%sp + 8]
"10000100011000100001000000000000",	-- 7527: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 7528: 	lw	%r2, [%r2 + 0]
"00111011110110110000000000000111",	-- 7529: 	lw	%r27, [%sp + 7]
"00111111111111100000000000001111",	-- 7530: 	sw	%ra, [%sp + 15]
"00111011011110100000000000000000",	-- 7531: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010000",	-- 7532: 	addi	%sp, %sp, 16
"01010011010000000000000000000000",	-- 7533: 	jalr	%r26
"10101011110111100000000000010000",	-- 7534: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 7535: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 7536: 	lli	%r2, 0
"00101000001000100000000000110100",	-- 7537: 	bneq	%r1, %r2, bneq_else.9183
"00111011110000010000000000001101",	-- 7538: 	lw	%r1, [%sp + 13]
"00111111111111100000000000001111",	-- 7539: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 7540: 	addi	%sp, %sp, 16
"01011000000000000000011010111010",	-- 7541: 	jal	d_vec.2683
"10101011110111100000000000010000",	-- 7542: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 7543: 	lw	%ra, [%sp + 15]
"10000100000000010001000000000000",	-- 7544: 	add	%r2, %r0, %r1
"00111011110000010000000000000110",	-- 7545: 	lw	%r1, [%sp + 6]
"00111111111111100000000000001111",	-- 7546: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 7547: 	addi	%sp, %sp, 16
"01011000000000000000010110100101",	-- 7548: 	jal	veciprod.2597
"10101011110111100000000000010000",	-- 7549: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 7550: 	lw	%ra, [%sp + 15]
"00111011110000010000000000001001",	-- 7551: 	lw	%r1, [%sp + 9]
"10110000000111100000000000001111",	-- 7552: 	sf	%f0, [%sp + 15]
"00111111111111100000000000010000",	-- 7553: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 7554: 	addi	%sp, %sp, 17
"01011000000000000000011011000010",	-- 7555: 	jal	r_bright.2691
"10101011110111100000000000010001",	-- 7556: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 7557: 	lw	%ra, [%sp + 16]
"10010011110000010000000000000101",	-- 7558: 	lf	%f1, [%sp + 5]
"11101000000000010001000000000000",	-- 7559: 	mulf	%f2, %f0, %f1
"10010011110000110000000000001111",	-- 7560: 	lf	%f3, [%sp + 15]
"11101000010000110001000000000000",	-- 7561: 	mulf	%f2, %f2, %f3
"00111011110000010000000000001101",	-- 7562: 	lw	%r1, [%sp + 13]
"10110000010111100000000000010000",	-- 7563: 	sf	%f2, [%sp + 16]
"10110000000111100000000000010001",	-- 7564: 	sf	%f0, [%sp + 17]
"00111111111111100000000000010010",	-- 7565: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 7566: 	addi	%sp, %sp, 19
"01011000000000000000011010111010",	-- 7567: 	jal	d_vec.2683
"10101011110111100000000000010011",	-- 7568: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 7569: 	lw	%ra, [%sp + 18]
"10000100000000010001000000000000",	-- 7570: 	add	%r2, %r0, %r1
"00111011110000010000000000000100",	-- 7571: 	lw	%r1, [%sp + 4]
"00111111111111100000000000010010",	-- 7572: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 7573: 	addi	%sp, %sp, 19
"01011000000000000000010110100101",	-- 7574: 	jal	veciprod.2597
"10101011110111100000000000010011",	-- 7575: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 7576: 	lw	%ra, [%sp + 18]
"10010011110000010000000000010001",	-- 7577: 	lf	%f1, [%sp + 17]
"11101000001000000000100000000000",	-- 7578: 	mulf	%f1, %f1, %f0
"10010011110000000000000000010000",	-- 7579: 	lf	%f0, [%sp + 16]
"10010011110000100000000000000010",	-- 7580: 	lf	%f2, [%sp + 2]
"00111011110110110000000000000011",	-- 7581: 	lw	%r27, [%sp + 3]
"00111111111111100000000000010010",	-- 7582: 	sw	%ra, [%sp + 18]
"00111011011110100000000000000000",	-- 7583: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010011",	-- 7584: 	addi	%sp, %sp, 19
"01010011010000000000000000000000",	-- 7585: 	jalr	%r26
"10101011110111100000000000010011",	-- 7586: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 7587: 	lw	%ra, [%sp + 18]
"01010100000000000001110110100101",	-- 7588: 	j	bneq_cont.9184
	-- bneq_else.9183:
	-- bneq_cont.9184:
"01010100000000000001110110100110",	-- 7589: 	j	bneq_cont.9182
	-- bneq_else.9181:
	-- bneq_cont.9182:
	-- bneq_cont.9180:
"11001100000000010000000000000001",	-- 7590: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 7591: 	lw	%r2, [%sp + 1]
"10001000010000010000100000000000",	-- 7592: 	sub	%r1, %r2, %r1
"10010011110000000000000000000101",	-- 7593: 	lf	%f0, [%sp + 5]
"10010011110000010000000000000010",	-- 7594: 	lf	%f1, [%sp + 2]
"00111011110000100000000000000100",	-- 7595: 	lw	%r2, [%sp + 4]
"00111011110110110000000000000000",	-- 7596: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 7597: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 7598: 	jr	%r26
	-- bgt_else.9178:
"01001111111000000000000000000000",	-- 7599: 	jr	%ra
	-- trace_ray.2903:
"00111011011001000000000000010100",	-- 7600: 	lw	%r4, [%r27 + 20]
"00111011011001010000000000010011",	-- 7601: 	lw	%r5, [%r27 + 19]
"00111011011001100000000000010010",	-- 7602: 	lw	%r6, [%r27 + 18]
"00111011011001110000000000010001",	-- 7603: 	lw	%r7, [%r27 + 17]
"00111011011010000000000000010000",	-- 7604: 	lw	%r8, [%r27 + 16]
"00111011011010010000000000001111",	-- 7605: 	lw	%r9, [%r27 + 15]
"00111011011010100000000000001110",	-- 7606: 	lw	%r10, [%r27 + 14]
"00111011011010110000000000001101",	-- 7607: 	lw	%r11, [%r27 + 13]
"00111011011011000000000000001100",	-- 7608: 	lw	%r12, [%r27 + 12]
"00111011011011010000000000001011",	-- 7609: 	lw	%r13, [%r27 + 11]
"00111011011011100000000000001010",	-- 7610: 	lw	%r14, [%r27 + 10]
"00111011011011110000000000001001",	-- 7611: 	lw	%r15, [%r27 + 9]
"00111011011100000000000000001000",	-- 7612: 	lw	%r16, [%r27 + 8]
"00111011011100010000000000000111",	-- 7613: 	lw	%r17, [%r27 + 7]
"00111011011100100000000000000110",	-- 7614: 	lw	%r18, [%r27 + 6]
"00111011011100110000000000000101",	-- 7615: 	lw	%r19, [%r27 + 5]
"00111011011101000000000000000100",	-- 7616: 	lw	%r20, [%r27 + 4]
"00111011011101010000000000000011",	-- 7617: 	lw	%r21, [%r27 + 3]
"00111011011101100000000000000010",	-- 7618: 	lw	%r22, [%r27 + 2]
"00111011011101110000000000000001",	-- 7619: 	lw	%r23, [%r27 + 1]
"11001100000110000000000000000100",	-- 7620: 	lli	%r24, 4
"00110000001110000000000110101111",	-- 7621: 	bgt	%r1, %r24, bgt_else.9186
"00111111011111100000000000000000",	-- 7622: 	sw	%r27, [%sp + 0]
"10110000001111100000000000000001",	-- 7623: 	sf	%f1, [%sp + 1]
"00111100110111100000000000000010",	-- 7624: 	sw	%r6, [%sp + 2]
"00111100101111100000000000000011",	-- 7625: 	sw	%r5, [%sp + 3]
"00111101111111100000000000000100",	-- 7626: 	sw	%r15, [%sp + 4]
"00111101010111100000000000000101",	-- 7627: 	sw	%r10, [%sp + 5]
"00111110111111100000000000000110",	-- 7628: 	sw	%r23, [%sp + 6]
"00111101001111100000000000000111",	-- 7629: 	sw	%r9, [%sp + 7]
"00111101100111100000000000001000",	-- 7630: 	sw	%r12, [%sp + 8]
"00111101110111100000000000001001",	-- 7631: 	sw	%r14, [%sp + 9]
"00111100111111100000000000001010",	-- 7632: 	sw	%r7, [%sp + 10]
"00111100011111100000000000001011",	-- 7633: 	sw	%r3, [%sp + 11]
"00111110010111100000000000001100",	-- 7634: 	sw	%r18, [%sp + 12]
"00111100100111100000000000001101",	-- 7635: 	sw	%r4, [%sp + 13]
"00111110011111100000000000001110",	-- 7636: 	sw	%r19, [%sp + 14]
"00111101000111100000000000001111",	-- 7637: 	sw	%r8, [%sp + 15]
"00111110101111100000000000010000",	-- 7638: 	sw	%r21, [%sp + 16]
"00111101101111100000000000010001",	-- 7639: 	sw	%r13, [%sp + 17]
"00111110100111100000000000010010",	-- 7640: 	sw	%r20, [%sp + 18]
"00111101011111100000000000010011",	-- 7641: 	sw	%r11, [%sp + 19]
"00111110110111100000000000010100",	-- 7642: 	sw	%r22, [%sp + 20]
"10110000000111100000000000010101",	-- 7643: 	sf	%f0, [%sp + 21]
"00111110000111100000000000010110",	-- 7644: 	sw	%r16, [%sp + 22]
"00111100001111100000000000010111",	-- 7645: 	sw	%r1, [%sp + 23]
"00111100010111100000000000011000",	-- 7646: 	sw	%r2, [%sp + 24]
"00111110001111100000000000011001",	-- 7647: 	sw	%r17, [%sp + 25]
"10000100000000110000100000000000",	-- 7648: 	add	%r1, %r0, %r3
"00111111111111100000000000011010",	-- 7649: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 7650: 	addi	%sp, %sp, 27
"01011000000000000000011010100110",	-- 7651: 	jal	p_surface_ids.2668
"10101011110111100000000000011011",	-- 7652: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 7653: 	lw	%ra, [%sp + 26]
"00111011110000100000000000011000",	-- 7654: 	lw	%r2, [%sp + 24]
"00111011110110110000000000011001",	-- 7655: 	lw	%r27, [%sp + 25]
"00111100001111100000000000011010",	-- 7656: 	sw	%r1, [%sp + 26]
"10000100000000100000100000000000",	-- 7657: 	add	%r1, %r0, %r2
"00111111111111100000000000011011",	-- 7658: 	sw	%ra, [%sp + 27]
"00111011011110100000000000000000",	-- 7659: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000011100",	-- 7660: 	addi	%sp, %sp, 28
"01010011010000000000000000000000",	-- 7661: 	jalr	%r26
"10101011110111100000000000011100",	-- 7662: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 7663: 	lw	%ra, [%sp + 27]
"11001100000000100000000000000000",	-- 7664: 	lli	%r2, 0
"00101000001000100000000001000101",	-- 7665: 	bneq	%r1, %r2, bneq_else.9187
"11001100000000011111111111111111",	-- 7666: 	lli	%r1, -1
"11001000000000011111111111111111",	-- 7667: 	lhi	%r1, -1
"00111011110000100000000000010111",	-- 7668: 	lw	%r2, [%sp + 23]
"00111011110000110000000000011010",	-- 7669: 	lw	%r3, [%sp + 26]
"10000100011000100001100000000000",	-- 7670: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 7671: 	sw	%r1, [%r3 + 0]
"11001100000000010000000000000000",	-- 7672: 	lli	%r1, 0
"00101000010000010000000000000010",	-- 7673: 	bneq	%r2, %r1, bneq_else.9188
"01001111111000000000000000000000",	-- 7674: 	jr	%ra
	-- bneq_else.9188:
"00111011110000010000000000011000",	-- 7675: 	lw	%r1, [%sp + 24]
"00111011110000100000000000010110",	-- 7676: 	lw	%r2, [%sp + 22]
"00111111111111100000000000011011",	-- 7677: 	sw	%ra, [%sp + 27]
"10100111110111100000000000011100",	-- 7678: 	addi	%sp, %sp, 28
"01011000000000000000010110100101",	-- 7679: 	jal	veciprod.2597
"10101011110111100000000000011100",	-- 7680: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 7681: 	lw	%ra, [%sp + 27]
"00111111111111100000000000011011",	-- 7682: 	sw	%ra, [%sp + 27]
"10100111110111100000000000011100",	-- 7683: 	addi	%sp, %sp, 28
"01011000000000000010101001001111",	-- 7684: 	jal	yj_fneg
"10101011110111100000000000011100",	-- 7685: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 7686: 	lw	%ra, [%sp + 27]
"10110000000111100000000000011011",	-- 7687: 	sf	%f0, [%sp + 27]
"00111111111111100000000000011100",	-- 7688: 	sw	%ra, [%sp + 28]
"10100111110111100000000000011101",	-- 7689: 	addi	%sp, %sp, 29
"01011000000000000000010011010100",	-- 7690: 	jal	fispos.2522
"10101011110111100000000000011101",	-- 7691: 	subi	%sp, %sp, 29
"00111011110111110000000000011100",	-- 7692: 	lw	%ra, [%sp + 28]
"11001100000000100000000000000000",	-- 7693: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 7694: 	bneq	%r1, %r2, bneq_else.9190
"01001111111000000000000000000000",	-- 7695: 	jr	%ra
	-- bneq_else.9190:
"10010011110000000000000000011011",	-- 7696: 	lf	%f0, [%sp + 27]
"00111111111111100000000000011100",	-- 7697: 	sw	%ra, [%sp + 28]
"10100111110111100000000000011101",	-- 7698: 	addi	%sp, %sp, 29
"01011000000000000000010011101111",	-- 7699: 	jal	fsqr.2530
"10101011110111100000000000011101",	-- 7700: 	subi	%sp, %sp, 29
"00111011110111110000000000011100",	-- 7701: 	lw	%ra, [%sp + 28]
"10010011110000010000000000011011",	-- 7702: 	lf	%f1, [%sp + 27]
"11101000000000010000000000000000",	-- 7703: 	mulf	%f0, %f0, %f1
"10010011110000010000000000010101",	-- 7704: 	lf	%f1, [%sp + 21]
"11101000000000010000000000000000",	-- 7705: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000000",	-- 7706: 	lli	%r1, 0
"00111011110000100000000000010100",	-- 7707: 	lw	%r2, [%sp + 20]
"10000100010000010000100000000000",	-- 7708: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 7709: 	lf	%f1, [%r1 + 0]
"11101000000000010000000000000000",	-- 7710: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000000",	-- 7711: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 7712: 	lli	%r2, 0
"00111011110000110000000000010011",	-- 7713: 	lw	%r3, [%sp + 19]
"10000100011000100001000000000000",	-- 7714: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 7715: 	lf	%f1, [%r2 + 0]
"11100000001000000000100000000000",	-- 7716: 	addf	%f1, %f1, %f0
"10000100011000010000100000000000",	-- 7717: 	add	%r1, %r3, %r1
"10110000001000010000000000000000",	-- 7718: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000001",	-- 7719: 	lli	%r1, 1
"11001100000000100000000000000001",	-- 7720: 	lli	%r2, 1
"10000100011000100001000000000000",	-- 7721: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 7722: 	lf	%f1, [%r2 + 0]
"11100000001000000000100000000000",	-- 7723: 	addf	%f1, %f1, %f0
"10000100011000010000100000000000",	-- 7724: 	add	%r1, %r3, %r1
"10110000001000010000000000000000",	-- 7725: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 7726: 	lli	%r1, 2
"11001100000000100000000000000010",	-- 7727: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 7728: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 7729: 	lf	%f1, [%r2 + 0]
"11100000001000000000000000000000",	-- 7730: 	addf	%f0, %f1, %f0
"10000100011000010000100000000000",	-- 7731: 	add	%r1, %r3, %r1
"10110000000000010000000000000000",	-- 7732: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 7733: 	jr	%ra
	-- bneq_else.9187:
"11001100000000010000000000000000",	-- 7734: 	lli	%r1, 0
"00111011110000100000000000010010",	-- 7735: 	lw	%r2, [%sp + 18]
"10000100010000010000100000000000",	-- 7736: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 7737: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000010001",	-- 7738: 	lw	%r2, [%sp + 17]
"10000100010000010001000000000000",	-- 7739: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 7740: 	lw	%r2, [%r2 + 0]
"00111100001111100000000000011100",	-- 7741: 	sw	%r1, [%sp + 28]
"00111100010111100000000000011101",	-- 7742: 	sw	%r2, [%sp + 29]
"10000100000000100000100000000000",	-- 7743: 	add	%r1, %r0, %r2
"00111111111111100000000000011110",	-- 7744: 	sw	%ra, [%sp + 30]
"10100111110111100000000000011111",	-- 7745: 	addi	%sp, %sp, 31
"01011000000000000000011001010010",	-- 7746: 	jal	o_reflectiontype.2626
"10101011110111100000000000011111",	-- 7747: 	subi	%sp, %sp, 31
"00111011110111110000000000011110",	-- 7748: 	lw	%ra, [%sp + 30]
"00111011110000100000000000011101",	-- 7749: 	lw	%r2, [%sp + 29]
"00111100001111100000000000011110",	-- 7750: 	sw	%r1, [%sp + 30]
"10000100000000100000100000000000",	-- 7751: 	add	%r1, %r0, %r2
"00111111111111100000000000011111",	-- 7752: 	sw	%ra, [%sp + 31]
"10100111110111100000000000100000",	-- 7753: 	addi	%sp, %sp, 32
"01011000000000000000011001111000",	-- 7754: 	jal	o_diffuse.2646
"10101011110111100000000000100000",	-- 7755: 	subi	%sp, %sp, 32
"00111011110111110000000000011111",	-- 7756: 	lw	%ra, [%sp + 31]
"10010011110000010000000000010101",	-- 7757: 	lf	%f1, [%sp + 21]
"11101000000000010000000000000000",	-- 7758: 	mulf	%f0, %f0, %f1
"00111011110000010000000000011101",	-- 7759: 	lw	%r1, [%sp + 29]
"00111011110000100000000000011000",	-- 7760: 	lw	%r2, [%sp + 24]
"00111011110110110000000000010000",	-- 7761: 	lw	%r27, [%sp + 16]
"10110000000111100000000000011111",	-- 7762: 	sf	%f0, [%sp + 31]
"00111111111111100000000000100000",	-- 7763: 	sw	%ra, [%sp + 32]
"00111011011110100000000000000000",	-- 7764: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100001",	-- 7765: 	addi	%sp, %sp, 33
"01010011010000000000000000000000",	-- 7766: 	jalr	%r26
"10101011110111100000000000100001",	-- 7767: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7768: 	lw	%ra, [%sp + 32]
"00111011110000010000000000001111",	-- 7769: 	lw	%r1, [%sp + 15]
"00111011110000100000000000001110",	-- 7770: 	lw	%r2, [%sp + 14]
"00111111111111100000000000100000",	-- 7771: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 7772: 	addi	%sp, %sp, 33
"01011000000000000000010100111011",	-- 7773: 	jal	veccpy.2586
"10101011110111100000000000100001",	-- 7774: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7775: 	lw	%ra, [%sp + 32]
"00111011110000010000000000011101",	-- 7776: 	lw	%r1, [%sp + 29]
"00111011110000100000000000001110",	-- 7777: 	lw	%r2, [%sp + 14]
"00111011110110110000000000001101",	-- 7778: 	lw	%r27, [%sp + 13]
"00111111111111100000000000100000",	-- 7779: 	sw	%ra, [%sp + 32]
"00111011011110100000000000000000",	-- 7780: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100001",	-- 7781: 	addi	%sp, %sp, 33
"01010011010000000000000000000000",	-- 7782: 	jalr	%r26
"10101011110111100000000000100001",	-- 7783: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7784: 	lw	%ra, [%sp + 32]
"11001100000000010000000000000100",	-- 7785: 	lli	%r1, 4
"00111011110000100000000000011100",	-- 7786: 	lw	%r2, [%sp + 28]
"10001100010000010000100000000000",	-- 7787: 	mul	%r1, %r2, %r1
"11001100000000100000000000000000",	-- 7788: 	lli	%r2, 0
"00111011110000110000000000001100",	-- 7789: 	lw	%r3, [%sp + 12]
"10000100011000100001000000000000",	-- 7790: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 7791: 	lw	%r2, [%r2 + 0]
"10000100001000100000100000000000",	-- 7792: 	add	%r1, %r1, %r2
"00111011110000100000000000010111",	-- 7793: 	lw	%r2, [%sp + 23]
"00111011110000110000000000011010",	-- 7794: 	lw	%r3, [%sp + 26]
"10000100011000100010000000000000",	-- 7795: 	add	%r4, %r3, %r2
"00111100001001000000000000000000",	-- 7796: 	sw	%r1, [%r4 + 0]
"00111011110000010000000000001011",	-- 7797: 	lw	%r1, [%sp + 11]
"00111111111111100000000000100000",	-- 7798: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 7799: 	addi	%sp, %sp, 33
"01011000000000000000011010100100",	-- 7800: 	jal	p_intersection_points.2666
"10101011110111100000000000100001",	-- 7801: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7802: 	lw	%ra, [%sp + 32]
"00111011110000100000000000010111",	-- 7803: 	lw	%r2, [%sp + 23]
"10000100001000100000100000000000",	-- 7804: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 7805: 	lw	%r1, [%r1 + 0]
"00111011110000110000000000001110",	-- 7806: 	lw	%r3, [%sp + 14]
"10000100000000110001000000000000",	-- 7807: 	add	%r2, %r0, %r3
"00111111111111100000000000100000",	-- 7808: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 7809: 	addi	%sp, %sp, 33
"01011000000000000000010100111011",	-- 7810: 	jal	veccpy.2586
"10101011110111100000000000100001",	-- 7811: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7812: 	lw	%ra, [%sp + 32]
"00111011110000010000000000001011",	-- 7813: 	lw	%r1, [%sp + 11]
"00111111111111100000000000100000",	-- 7814: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 7815: 	addi	%sp, %sp, 33
"01011000000000000000011010101000",	-- 7816: 	jal	p_calc_diffuse.2670
"10101011110111100000000000100001",	-- 7817: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7818: 	lw	%ra, [%sp + 32]
"00111011110000100000000000011101",	-- 7819: 	lw	%r2, [%sp + 29]
"00111100001111100000000000100000",	-- 7820: 	sw	%r1, [%sp + 32]
"10000100000000100000100000000000",	-- 7821: 	add	%r1, %r0, %r2
"00111111111111100000000000100001",	-- 7822: 	sw	%ra, [%sp + 33]
"10100111110111100000000000100010",	-- 7823: 	addi	%sp, %sp, 34
"01011000000000000000011001111000",	-- 7824: 	jal	o_diffuse.2646
"10101011110111100000000000100010",	-- 7825: 	subi	%sp, %sp, 34
"00111011110111110000000000100001",	-- 7826: 	lw	%ra, [%sp + 33]
"00010100000000010000000000000000",	-- 7827: 	llif	%f1, 0.500000
"00010000000000010011111100000000",	-- 7828: 	lhif	%f1, 0.500000
"00111111111111100000000000100001",	-- 7829: 	sw	%ra, [%sp + 33]
"10100111110111100000000000100010",	-- 7830: 	addi	%sp, %sp, 34
"01011000000000000000010011110001",	-- 7831: 	jal	fless.2532
"10101011110111100000000000100010",	-- 7832: 	subi	%sp, %sp, 34
"00111011110111110000000000100001",	-- 7833: 	lw	%ra, [%sp + 33]
"11001100000000100000000000000000",	-- 7834: 	lli	%r2, 0
"00101000001000100000000000110111",	-- 7835: 	bneq	%r1, %r2, bneq_else.9193
"11001100000000010000000000000001",	-- 7836: 	lli	%r1, 1
"00111011110000100000000000010111",	-- 7837: 	lw	%r2, [%sp + 23]
"00111011110000110000000000100000",	-- 7838: 	lw	%r3, [%sp + 32]
"10000100011000100001100000000000",	-- 7839: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 7840: 	sw	%r1, [%r3 + 0]
"00111011110000010000000000001011",	-- 7841: 	lw	%r1, [%sp + 11]
"00111111111111100000000000100001",	-- 7842: 	sw	%ra, [%sp + 33]
"10100111110111100000000000100010",	-- 7843: 	addi	%sp, %sp, 34
"01011000000000000000011010101010",	-- 7844: 	jal	p_energy.2672
"10101011110111100000000000100010",	-- 7845: 	subi	%sp, %sp, 34
"00111011110111110000000000100001",	-- 7846: 	lw	%ra, [%sp + 33]
"00111011110000100000000000010111",	-- 7847: 	lw	%r2, [%sp + 23]
"10000100001000100001100000000000",	-- 7848: 	add	%r3, %r1, %r2
"00111000011000110000000000000000",	-- 7849: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000001010",	-- 7850: 	lw	%r4, [%sp + 10]
"00111100001111100000000000100001",	-- 7851: 	sw	%r1, [%sp + 33]
"10000100000001000001000000000000",	-- 7852: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 7853: 	add	%r1, %r0, %r3
"00111111111111100000000000100010",	-- 7854: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 7855: 	addi	%sp, %sp, 35
"01011000000000000000010100111011",	-- 7856: 	jal	veccpy.2586
"10101011110111100000000000100011",	-- 7857: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 7858: 	lw	%ra, [%sp + 34]
"00111011110000010000000000010111",	-- 7859: 	lw	%r1, [%sp + 23]
"00111011110000100000000000100001",	-- 7860: 	lw	%r2, [%sp + 33]
"10000100010000010001000000000000",	-- 7861: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 7862: 	lw	%r2, [%r2 + 0]
"00010100000000001111101111001110",	-- 7863: 	llif	%f0, 0.003906
"00010000000000000011101101111111",	-- 7864: 	lhif	%f0, 0.003906
"10010011110000010000000000011111",	-- 7865: 	lf	%f1, [%sp + 31]
"11101000000000010000000000000000",	-- 7866: 	mulf	%f0, %f0, %f1
"10000100000000100000100000000000",	-- 7867: 	add	%r1, %r0, %r2
"00111111111111100000000000100010",	-- 7868: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 7869: 	addi	%sp, %sp, 35
"01011000000000000000011000001101",	-- 7870: 	jal	vecscale.2615
"10101011110111100000000000100011",	-- 7871: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 7872: 	lw	%ra, [%sp + 34]
"00111011110000010000000000001011",	-- 7873: 	lw	%r1, [%sp + 11]
"00111111111111100000000000100010",	-- 7874: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 7875: 	addi	%sp, %sp, 35
"01011000000000000000011010111000",	-- 7876: 	jal	p_nvectors.2681
"10101011110111100000000000100011",	-- 7877: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 7878: 	lw	%ra, [%sp + 34]
"00111011110000100000000000010111",	-- 7879: 	lw	%r2, [%sp + 23]
"10000100001000100000100000000000",	-- 7880: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 7881: 	lw	%r1, [%r1 + 0]
"00111011110000110000000000001001",	-- 7882: 	lw	%r3, [%sp + 9]
"10000100000000110001000000000000",	-- 7883: 	add	%r2, %r0, %r3
"00111111111111100000000000100010",	-- 7884: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 7885: 	addi	%sp, %sp, 35
"01011000000000000000010100111011",	-- 7886: 	jal	veccpy.2586
"10101011110111100000000000100011",	-- 7887: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 7888: 	lw	%ra, [%sp + 34]
"01010100000000000001111011010111",	-- 7889: 	j	bneq_cont.9194
	-- bneq_else.9193:
"11001100000000010000000000000000",	-- 7890: 	lli	%r1, 0
"00111011110000100000000000010111",	-- 7891: 	lw	%r2, [%sp + 23]
"00111011110000110000000000100000",	-- 7892: 	lw	%r3, [%sp + 32]
"10000100011000100001100000000000",	-- 7893: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 7894: 	sw	%r1, [%r3 + 0]
	-- bneq_cont.9194:
"00010100000000000000000000000000",	-- 7895: 	llif	%f0, -2.000000
"00010000000000001100000000000000",	-- 7896: 	lhif	%f0, -2.000000
"00111011110000010000000000011000",	-- 7897: 	lw	%r1, [%sp + 24]
"00111011110000100000000000001001",	-- 7898: 	lw	%r2, [%sp + 9]
"10110000000111100000000000100010",	-- 7899: 	sf	%f0, [%sp + 34]
"00111111111111100000000000100011",	-- 7900: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 7901: 	addi	%sp, %sp, 36
"01011000000000000000010110100101",	-- 7902: 	jal	veciprod.2597
"10101011110111100000000000100100",	-- 7903: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 7904: 	lw	%ra, [%sp + 35]
"10010011110000010000000000100010",	-- 7905: 	lf	%f1, [%sp + 34]
"11101000001000000000000000000000",	-- 7906: 	mulf	%f0, %f1, %f0
"00111011110000010000000000011000",	-- 7907: 	lw	%r1, [%sp + 24]
"00111011110000100000000000001001",	-- 7908: 	lw	%r2, [%sp + 9]
"00111111111111100000000000100011",	-- 7909: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 7910: 	addi	%sp, %sp, 36
"01011000000000000000010111001100",	-- 7911: 	jal	vecaccum.2605
"10101011110111100000000000100100",	-- 7912: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 7913: 	lw	%ra, [%sp + 35]
"00111011110000010000000000011101",	-- 7914: 	lw	%r1, [%sp + 29]
"00111111111111100000000000100011",	-- 7915: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 7916: 	addi	%sp, %sp, 36
"01011000000000000000011001111101",	-- 7917: 	jal	o_hilight.2648
"10101011110111100000000000100100",	-- 7918: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 7919: 	lw	%ra, [%sp + 35]
"10010011110000010000000000010101",	-- 7920: 	lf	%f1, [%sp + 21]
"11101000001000000000000000000000",	-- 7921: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 7922: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 7923: 	lli	%r2, 0
"00111011110000110000000000001000",	-- 7924: 	lw	%r3, [%sp + 8]
"10000100011000100001000000000000",	-- 7925: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 7926: 	lw	%r2, [%r2 + 0]
"00111011110110110000000000000111",	-- 7927: 	lw	%r27, [%sp + 7]
"10110000000111100000000000100011",	-- 7928: 	sf	%f0, [%sp + 35]
"00111111111111100000000000100100",	-- 7929: 	sw	%ra, [%sp + 36]
"00111011011110100000000000000000",	-- 7930: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100101",	-- 7931: 	addi	%sp, %sp, 37
"01010011010000000000000000000000",	-- 7932: 	jalr	%r26
"10101011110111100000000000100101",	-- 7933: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 7934: 	lw	%ra, [%sp + 36]
"11001100000000100000000000000000",	-- 7935: 	lli	%r2, 0
"00101000001000100000000000100111",	-- 7936: 	bneq	%r1, %r2, bneq_else.9195
"00111011110000010000000000001001",	-- 7937: 	lw	%r1, [%sp + 9]
"00111011110000100000000000010110",	-- 7938: 	lw	%r2, [%sp + 22]
"00111111111111100000000000100100",	-- 7939: 	sw	%ra, [%sp + 36]
"10100111110111100000000000100101",	-- 7940: 	addi	%sp, %sp, 37
"01011000000000000000010110100101",	-- 7941: 	jal	veciprod.2597
"10101011110111100000000000100101",	-- 7942: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 7943: 	lw	%ra, [%sp + 36]
"00111111111111100000000000100100",	-- 7944: 	sw	%ra, [%sp + 36]
"10100111110111100000000000100101",	-- 7945: 	addi	%sp, %sp, 37
"01011000000000000010101001001111",	-- 7946: 	jal	yj_fneg
"10101011110111100000000000100101",	-- 7947: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 7948: 	lw	%ra, [%sp + 36]
"10010011110000010000000000011111",	-- 7949: 	lf	%f1, [%sp + 31]
"11101000000000010000000000000000",	-- 7950: 	mulf	%f0, %f0, %f1
"00111011110000010000000000011000",	-- 7951: 	lw	%r1, [%sp + 24]
"00111011110000100000000000010110",	-- 7952: 	lw	%r2, [%sp + 22]
"10110000000111100000000000100100",	-- 7953: 	sf	%f0, [%sp + 36]
"00111111111111100000000000100101",	-- 7954: 	sw	%ra, [%sp + 37]
"10100111110111100000000000100110",	-- 7955: 	addi	%sp, %sp, 38
"01011000000000000000010110100101",	-- 7956: 	jal	veciprod.2597
"10101011110111100000000000100110",	-- 7957: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 7958: 	lw	%ra, [%sp + 37]
"00111111111111100000000000100101",	-- 7959: 	sw	%ra, [%sp + 37]
"10100111110111100000000000100110",	-- 7960: 	addi	%sp, %sp, 38
"01011000000000000010101001001111",	-- 7961: 	jal	yj_fneg
"10101011110111100000000000100110",	-- 7962: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 7963: 	lw	%ra, [%sp + 37]
"00001100000000010000000000000000",	-- 7964: 	movf	%f1, %f0
"10010011110000000000000000100100",	-- 7965: 	lf	%f0, [%sp + 36]
"10010011110000100000000000100011",	-- 7966: 	lf	%f2, [%sp + 35]
"00111011110110110000000000000110",	-- 7967: 	lw	%r27, [%sp + 6]
"00111111111111100000000000100101",	-- 7968: 	sw	%ra, [%sp + 37]
"00111011011110100000000000000000",	-- 7969: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100110",	-- 7970: 	addi	%sp, %sp, 38
"01010011010000000000000000000000",	-- 7971: 	jalr	%r26
"10101011110111100000000000100110",	-- 7972: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 7973: 	lw	%ra, [%sp + 37]
"01010100000000000001111100100111",	-- 7974: 	j	bneq_cont.9196
	-- bneq_else.9195:
	-- bneq_cont.9196:
"00111011110000010000000000001110",	-- 7975: 	lw	%r1, [%sp + 14]
"00111011110110110000000000000101",	-- 7976: 	lw	%r27, [%sp + 5]
"00111111111111100000000000100101",	-- 7977: 	sw	%ra, [%sp + 37]
"00111011011110100000000000000000",	-- 7978: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100110",	-- 7979: 	addi	%sp, %sp, 38
"01010011010000000000000000000000",	-- 7980: 	jalr	%r26
"10101011110111100000000000100110",	-- 7981: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 7982: 	lw	%ra, [%sp + 37]
"11001100000000010000000000000000",	-- 7983: 	lli	%r1, 0
"00111011110000100000000000000100",	-- 7984: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 7985: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 7986: 	lw	%r1, [%r1 + 0]
"11001100000000100000000000000001",	-- 7987: 	lli	%r2, 1
"10001000001000100000100000000000",	-- 7988: 	sub	%r1, %r1, %r2
"10010011110000000000000000011111",	-- 7989: 	lf	%f0, [%sp + 31]
"10010011110000010000000000100011",	-- 7990: 	lf	%f1, [%sp + 35]
"00111011110000100000000000011000",	-- 7991: 	lw	%r2, [%sp + 24]
"00111011110110110000000000000011",	-- 7992: 	lw	%r27, [%sp + 3]
"00111111111111100000000000100101",	-- 7993: 	sw	%ra, [%sp + 37]
"00111011011110100000000000000000",	-- 7994: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100110",	-- 7995: 	addi	%sp, %sp, 38
"01010011010000000000000000000000",	-- 7996: 	jalr	%r26
"10101011110111100000000000100110",	-- 7997: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 7998: 	lw	%ra, [%sp + 37]
"00010100000000001100110011001101",	-- 7999: 	llif	%f0, 0.100000
"00010000000000000011110111001100",	-- 8000: 	lhif	%f0, 0.100000
"10010011110000010000000000010101",	-- 8001: 	lf	%f1, [%sp + 21]
"00111111111111100000000000100101",	-- 8002: 	sw	%ra, [%sp + 37]
"10100111110111100000000000100110",	-- 8003: 	addi	%sp, %sp, 38
"01011000000000000000010011110001",	-- 8004: 	jal	fless.2532
"10101011110111100000000000100110",	-- 8005: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 8006: 	lw	%ra, [%sp + 37]
"11001100000000100000000000000000",	-- 8007: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 8008: 	bneq	%r1, %r2, bneq_else.9197
"01001111111000000000000000000000",	-- 8009: 	jr	%ra
	-- bneq_else.9197:
"11001100000000010000000000000100",	-- 8010: 	lli	%r1, 4
"00111011110000100000000000010111",	-- 8011: 	lw	%r2, [%sp + 23]
"00110000001000100000000000000010",	-- 8012: 	bgt	%r1, %r2, bgt_else.9199
"01010100000000000001111101010101",	-- 8013: 	j	bgt_cont.9200
	-- bgt_else.9199:
"11001100000000010000000000000001",	-- 8014: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 8015: 	add	%r1, %r2, %r1
"11001100000000111111111111111111",	-- 8016: 	lli	%r3, -1
"11001000000000111111111111111111",	-- 8017: 	lhi	%r3, -1
"00111011110001000000000000011010",	-- 8018: 	lw	%r4, [%sp + 26]
"10000100100000010000100000000000",	-- 8019: 	add	%r1, %r4, %r1
"00111100011000010000000000000000",	-- 8020: 	sw	%r3, [%r1 + 0]
	-- bgt_cont.9200:
"11001100000000010000000000000010",	-- 8021: 	lli	%r1, 2
"00111011110000110000000000011110",	-- 8022: 	lw	%r3, [%sp + 30]
"00101000011000010000000000011100",	-- 8023: 	bneq	%r3, %r1, bneq_else.9201
"00010100000000000000000000000000",	-- 8024: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 8025: 	lhif	%f0, 1.000000
"00111011110000010000000000011101",	-- 8026: 	lw	%r1, [%sp + 29]
"10110000000111100000000000100101",	-- 8027: 	sf	%f0, [%sp + 37]
"00111111111111100000000000100110",	-- 8028: 	sw	%ra, [%sp + 38]
"10100111110111100000000000100111",	-- 8029: 	addi	%sp, %sp, 39
"01011000000000000000011001111000",	-- 8030: 	jal	o_diffuse.2646
"10101011110111100000000000100111",	-- 8031: 	subi	%sp, %sp, 39
"00111011110111110000000000100110",	-- 8032: 	lw	%ra, [%sp + 38]
"10010011110000010000000000100101",	-- 8033: 	lf	%f1, [%sp + 37]
"11100100001000000000000000000000",	-- 8034: 	subf	%f0, %f1, %f0
"10010011110000010000000000010101",	-- 8035: 	lf	%f1, [%sp + 21]
"11101000001000000000000000000000",	-- 8036: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 8037: 	lli	%r1, 1
"00111011110000100000000000010111",	-- 8038: 	lw	%r2, [%sp + 23]
"10000100010000010000100000000000",	-- 8039: 	add	%r1, %r2, %r1
"11001100000000100000000000000000",	-- 8040: 	lli	%r2, 0
"00111011110000110000000000000010",	-- 8041: 	lw	%r3, [%sp + 2]
"10000100011000100001000000000000",	-- 8042: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 8043: 	lf	%f1, [%r2 + 0]
"10010011110000100000000000000001",	-- 8044: 	lf	%f2, [%sp + 1]
"11100000010000010000100000000000",	-- 8045: 	addf	%f1, %f2, %f1
"00111011110000100000000000011000",	-- 8046: 	lw	%r2, [%sp + 24]
"00111011110000110000000000001011",	-- 8047: 	lw	%r3, [%sp + 11]
"00111011110110110000000000000000",	-- 8048: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 8049: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8050: 	jr	%r26
	-- bneq_else.9201:
"01001111111000000000000000000000",	-- 8051: 	jr	%ra
	-- bgt_else.9186:
"01001111111000000000000000000000",	-- 8052: 	jr	%ra
	-- trace_diffuse_ray.2909:
"00111011011000100000000000001100",	-- 8053: 	lw	%r2, [%r27 + 12]
"00111011011000110000000000001011",	-- 8054: 	lw	%r3, [%r27 + 11]
"00111011011001000000000000001010",	-- 8055: 	lw	%r4, [%r27 + 10]
"00111011011001010000000000001001",	-- 8056: 	lw	%r5, [%r27 + 9]
"00111011011001100000000000001000",	-- 8057: 	lw	%r6, [%r27 + 8]
"00111011011001110000000000000111",	-- 8058: 	lw	%r7, [%r27 + 7]
"00111011011010000000000000000110",	-- 8059: 	lw	%r8, [%r27 + 6]
"00111011011010010000000000000101",	-- 8060: 	lw	%r9, [%r27 + 5]
"00111011011010100000000000000100",	-- 8061: 	lw	%r10, [%r27 + 4]
"00111011011010110000000000000011",	-- 8062: 	lw	%r11, [%r27 + 3]
"00111011011011000000000000000010",	-- 8063: 	lw	%r12, [%r27 + 2]
"00111011011011010000000000000001",	-- 8064: 	lw	%r13, [%r27 + 1]
"00111100011111100000000000000000",	-- 8065: 	sw	%r3, [%sp + 0]
"00111101101111100000000000000001",	-- 8066: 	sw	%r13, [%sp + 1]
"10110000000111100000000000000010",	-- 8067: 	sf	%f0, [%sp + 2]
"00111101000111100000000000000011",	-- 8068: 	sw	%r8, [%sp + 3]
"00111100111111100000000000000100",	-- 8069: 	sw	%r7, [%sp + 4]
"00111100100111100000000000000101",	-- 8070: 	sw	%r4, [%sp + 5]
"00111100101111100000000000000110",	-- 8071: 	sw	%r5, [%sp + 6]
"00111101010111100000000000000111",	-- 8072: 	sw	%r10, [%sp + 7]
"00111100010111100000000000001000",	-- 8073: 	sw	%r2, [%sp + 8]
"00111101100111100000000000001001",	-- 8074: 	sw	%r12, [%sp + 9]
"00111100001111100000000000001010",	-- 8075: 	sw	%r1, [%sp + 10]
"00111100110111100000000000001011",	-- 8076: 	sw	%r6, [%sp + 11]
"00111101011111100000000000001100",	-- 8077: 	sw	%r11, [%sp + 12]
"10000100000010011101100000000000",	-- 8078: 	add	%r27, %r0, %r9
"00111111111111100000000000001101",	-- 8079: 	sw	%ra, [%sp + 13]
"00111011011110100000000000000000",	-- 8080: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001110",	-- 8081: 	addi	%sp, %sp, 14
"01010011010000000000000000000000",	-- 8082: 	jalr	%r26
"10101011110111100000000000001110",	-- 8083: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 8084: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 8085: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 8086: 	bneq	%r1, %r2, bneq_else.9204
"01001111111000000000000000000000",	-- 8087: 	jr	%ra
	-- bneq_else.9204:
"11001100000000010000000000000000",	-- 8088: 	lli	%r1, 0
"00111011110000100000000000001100",	-- 8089: 	lw	%r2, [%sp + 12]
"10000100010000010000100000000000",	-- 8090: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8091: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000001011",	-- 8092: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 8093: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8094: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000001010",	-- 8095: 	lw	%r2, [%sp + 10]
"00111100001111100000000000001101",	-- 8096: 	sw	%r1, [%sp + 13]
"10000100000000100000100000000000",	-- 8097: 	add	%r1, %r0, %r2
"00111111111111100000000000001110",	-- 8098: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 8099: 	addi	%sp, %sp, 15
"01011000000000000000011010111010",	-- 8100: 	jal	d_vec.2683
"10101011110111100000000000001111",	-- 8101: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 8102: 	lw	%ra, [%sp + 14]
"10000100000000010001000000000000",	-- 8103: 	add	%r2, %r0, %r1
"00111011110000010000000000001101",	-- 8104: 	lw	%r1, [%sp + 13]
"00111011110110110000000000001001",	-- 8105: 	lw	%r27, [%sp + 9]
"00111111111111100000000000001110",	-- 8106: 	sw	%ra, [%sp + 14]
"00111011011110100000000000000000",	-- 8107: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001111",	-- 8108: 	addi	%sp, %sp, 15
"01010011010000000000000000000000",	-- 8109: 	jalr	%r26
"10101011110111100000000000001111",	-- 8110: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 8111: 	lw	%ra, [%sp + 14]
"00111011110000010000000000001101",	-- 8112: 	lw	%r1, [%sp + 13]
"00111011110000100000000000000111",	-- 8113: 	lw	%r2, [%sp + 7]
"00111011110110110000000000001000",	-- 8114: 	lw	%r27, [%sp + 8]
"00111111111111100000000000001110",	-- 8115: 	sw	%ra, [%sp + 14]
"00111011011110100000000000000000",	-- 8116: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001111",	-- 8117: 	addi	%sp, %sp, 15
"01010011010000000000000000000000",	-- 8118: 	jalr	%r26
"10101011110111100000000000001111",	-- 8119: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 8120: 	lw	%ra, [%sp + 14]
"11001100000000010000000000000000",	-- 8121: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 8122: 	lli	%r2, 0
"00111011110000110000000000000110",	-- 8123: 	lw	%r3, [%sp + 6]
"10000100011000100001000000000000",	-- 8124: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 8125: 	lw	%r2, [%r2 + 0]
"00111011110110110000000000000101",	-- 8126: 	lw	%r27, [%sp + 5]
"00111111111111100000000000001110",	-- 8127: 	sw	%ra, [%sp + 14]
"00111011011110100000000000000000",	-- 8128: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001111",	-- 8129: 	addi	%sp, %sp, 15
"01010011010000000000000000000000",	-- 8130: 	jalr	%r26
"10101011110111100000000000001111",	-- 8131: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 8132: 	lw	%ra, [%sp + 14]
"11001100000000100000000000000000",	-- 8133: 	lli	%r2, 0
"00101000001000100000000000100111",	-- 8134: 	bneq	%r1, %r2, bneq_else.9206
"00111011110000010000000000000100",	-- 8135: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000011",	-- 8136: 	lw	%r2, [%sp + 3]
"00111111111111100000000000001110",	-- 8137: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 8138: 	addi	%sp, %sp, 15
"01011000000000000000010110100101",	-- 8139: 	jal	veciprod.2597
"10101011110111100000000000001111",	-- 8140: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 8141: 	lw	%ra, [%sp + 14]
"00111111111111100000000000001110",	-- 8142: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 8143: 	addi	%sp, %sp, 15
"01011000000000000010101001001111",	-- 8144: 	jal	yj_fneg
"10101011110111100000000000001111",	-- 8145: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 8146: 	lw	%ra, [%sp + 14]
"10110000000111100000000000001110",	-- 8147: 	sf	%f0, [%sp + 14]
"00111111111111100000000000001111",	-- 8148: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 8149: 	addi	%sp, %sp, 16
"01011000000000000000010011010100",	-- 8150: 	jal	fispos.2522
"10101011110111100000000000010000",	-- 8151: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 8152: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 8153: 	lli	%r2, 0
"00101000001000100000000000000100",	-- 8154: 	bneq	%r1, %r2, bneq_else.9207
"00010100000000000000000000000000",	-- 8155: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 8156: 	lhif	%f0, 0.000000
"01010100000000000001111111011111",	-- 8157: 	j	bneq_cont.9208
	-- bneq_else.9207:
"10010011110000000000000000001110",	-- 8158: 	lf	%f0, [%sp + 14]
	-- bneq_cont.9208:
"10010011110000010000000000000010",	-- 8159: 	lf	%f1, [%sp + 2]
"11101000001000000000000000000000",	-- 8160: 	mulf	%f0, %f1, %f0
"00111011110000010000000000001101",	-- 8161: 	lw	%r1, [%sp + 13]
"10110000000111100000000000001111",	-- 8162: 	sf	%f0, [%sp + 15]
"00111111111111100000000000010000",	-- 8163: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 8164: 	addi	%sp, %sp, 17
"01011000000000000000011001111000",	-- 8165: 	jal	o_diffuse.2646
"10101011110111100000000000010001",	-- 8166: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 8167: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001111",	-- 8168: 	lf	%f1, [%sp + 15]
"11101000001000000000000000000000",	-- 8169: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 8170: 	lw	%r1, [%sp + 1]
"00111011110000100000000000000000",	-- 8171: 	lw	%r2, [%sp + 0]
"01010100000000000000010111001100",	-- 8172: 	j	vecaccum.2605
	-- bneq_else.9206:
"01001111111000000000000000000000",	-- 8173: 	jr	%ra
	-- iter_trace_diffuse_rays.2912:
"00111011011001010000000000000001",	-- 8174: 	lw	%r5, [%r27 + 1]
"11001100000001100000000000000000",	-- 8175: 	lli	%r6, 0
"00110000110001000000000001001000",	-- 8176: 	bgt	%r6, %r4, bgt_else.9210
"10000100001001000011000000000000",	-- 8177: 	add	%r6, %r1, %r4
"00111000110001100000000000000000",	-- 8178: 	lw	%r6, [%r6 + 0]
"00111100011111100000000000000000",	-- 8179: 	sw	%r3, [%sp + 0]
"00111111011111100000000000000001",	-- 8180: 	sw	%r27, [%sp + 1]
"00111100101111100000000000000010",	-- 8181: 	sw	%r5, [%sp + 2]
"00111100100111100000000000000011",	-- 8182: 	sw	%r4, [%sp + 3]
"00111100001111100000000000000100",	-- 8183: 	sw	%r1, [%sp + 4]
"00111100010111100000000000000101",	-- 8184: 	sw	%r2, [%sp + 5]
"10000100000001100000100000000000",	-- 8185: 	add	%r1, %r0, %r6
"00111111111111100000000000000110",	-- 8186: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8187: 	addi	%sp, %sp, 7
"01011000000000000000011010111010",	-- 8188: 	jal	d_vec.2683
"10101011110111100000000000000111",	-- 8189: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8190: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000101",	-- 8191: 	lw	%r2, [%sp + 5]
"00111111111111100000000000000110",	-- 8192: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8193: 	addi	%sp, %sp, 7
"01011000000000000000010110100101",	-- 8194: 	jal	veciprod.2597
"10101011110111100000000000000111",	-- 8195: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8196: 	lw	%ra, [%sp + 6]
"10110000000111100000000000000110",	-- 8197: 	sf	%f0, [%sp + 6]
"00111111111111100000000000000111",	-- 8198: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 8199: 	addi	%sp, %sp, 8
"01011000000000000000010011011011",	-- 8200: 	jal	fisneg.2524
"10101011110111100000000000001000",	-- 8201: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8202: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000000",	-- 8203: 	lli	%r2, 0
"00101000001000100000000000010010",	-- 8204: 	bneq	%r1, %r2, bneq_else.9211
"00111011110000010000000000000011",	-- 8205: 	lw	%r1, [%sp + 3]
"00111011110000100000000000000100",	-- 8206: 	lw	%r2, [%sp + 4]
"10000100010000010001100000000000",	-- 8207: 	add	%r3, %r2, %r1
"00111000011000110000000000000000",	-- 8208: 	lw	%r3, [%r3 + 0]
"00010100000000000000000000000000",	-- 8209: 	llif	%f0, 150.000000
"00010000000000000100001100010110",	-- 8210: 	lhif	%f0, 150.000000
"10010011110000010000000000000110",	-- 8211: 	lf	%f1, [%sp + 6]
"11101100001000000000000000000000",	-- 8212: 	divf	%f0, %f1, %f0
"00111011110110110000000000000010",	-- 8213: 	lw	%r27, [%sp + 2]
"10000100000000110000100000000000",	-- 8214: 	add	%r1, %r0, %r3
"00111111111111100000000000000111",	-- 8215: 	sw	%ra, [%sp + 7]
"00111011011110100000000000000000",	-- 8216: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001000",	-- 8217: 	addi	%sp, %sp, 8
"01010011010000000000000000000000",	-- 8218: 	jalr	%r26
"10101011110111100000000000001000",	-- 8219: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8220: 	lw	%ra, [%sp + 7]
"01010100000000000010000000101111",	-- 8221: 	j	bneq_cont.9212
	-- bneq_else.9211:
"11001100000000010000000000000001",	-- 8222: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 8223: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 8224: 	add	%r1, %r2, %r1
"00111011110000110000000000000100",	-- 8225: 	lw	%r3, [%sp + 4]
"10000100011000010000100000000000",	-- 8226: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 8227: 	lw	%r1, [%r1 + 0]
"00010100000000000000000000000000",	-- 8228: 	llif	%f0, -150.000000
"00010000000000001100001100010110",	-- 8229: 	lhif	%f0, -150.000000
"10010011110000010000000000000110",	-- 8230: 	lf	%f1, [%sp + 6]
"11101100001000000000000000000000",	-- 8231: 	divf	%f0, %f1, %f0
"00111011110110110000000000000010",	-- 8232: 	lw	%r27, [%sp + 2]
"00111111111111100000000000000111",	-- 8233: 	sw	%ra, [%sp + 7]
"00111011011110100000000000000000",	-- 8234: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001000",	-- 8235: 	addi	%sp, %sp, 8
"01010011010000000000000000000000",	-- 8236: 	jalr	%r26
"10101011110111100000000000001000",	-- 8237: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8238: 	lw	%ra, [%sp + 7]
	-- bneq_cont.9212:
"11001100000000010000000000000010",	-- 8239: 	lli	%r1, 2
"00111011110000100000000000000011",	-- 8240: 	lw	%r2, [%sp + 3]
"10001000010000010010000000000000",	-- 8241: 	sub	%r4, %r2, %r1
"00111011110000010000000000000100",	-- 8242: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000101",	-- 8243: 	lw	%r2, [%sp + 5]
"00111011110000110000000000000000",	-- 8244: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000001",	-- 8245: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 8246: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8247: 	jr	%r26
	-- bgt_else.9210:
"01001111111000000000000000000000",	-- 8248: 	jr	%ra
	-- trace_diffuse_rays.2917:
"00111011011001000000000000000010",	-- 8249: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 8250: 	lw	%r5, [%r27 + 1]
"00111100011111100000000000000000",	-- 8251: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 8252: 	sw	%r2, [%sp + 1]
"00111100001111100000000000000010",	-- 8253: 	sw	%r1, [%sp + 2]
"00111100101111100000000000000011",	-- 8254: 	sw	%r5, [%sp + 3]
"10000100000000110000100000000000",	-- 8255: 	add	%r1, %r0, %r3
"10000100000001001101100000000000",	-- 8256: 	add	%r27, %r0, %r4
"00111111111111100000000000000100",	-- 8257: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 8258: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 8259: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 8260: 	jalr	%r26
"10101011110111100000000000000101",	-- 8261: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 8262: 	lw	%ra, [%sp + 4]
"11001100000001000000000001110110",	-- 8263: 	lli	%r4, 118
"00111011110000010000000000000010",	-- 8264: 	lw	%r1, [%sp + 2]
"00111011110000100000000000000001",	-- 8265: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 8266: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000011",	-- 8267: 	lw	%r27, [%sp + 3]
"00111011011110100000000000000000",	-- 8268: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8269: 	jr	%r26
	-- trace_diffuse_ray_80percent.2921:
"00111011011001000000000000000010",	-- 8270: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 8271: 	lw	%r5, [%r27 + 1]
"11001100000001100000000000000000",	-- 8272: 	lli	%r6, 0
"00111100011111100000000000000000",	-- 8273: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 8274: 	sw	%r2, [%sp + 1]
"00111100100111100000000000000010",	-- 8275: 	sw	%r4, [%sp + 2]
"00111100101111100000000000000011",	-- 8276: 	sw	%r5, [%sp + 3]
"00111100001111100000000000000100",	-- 8277: 	sw	%r1, [%sp + 4]
"00101000001001100000000000000010",	-- 8278: 	bneq	%r1, %r6, bneq_else.9214
"01010100000000000010000001100011",	-- 8279: 	j	bneq_cont.9215
	-- bneq_else.9214:
"11001100000001100000000000000000",	-- 8280: 	lli	%r6, 0
"10000100101001100011000000000000",	-- 8281: 	add	%r6, %r5, %r6
"00111000110001100000000000000000",	-- 8282: 	lw	%r6, [%r6 + 0]
"10000100000001100000100000000000",	-- 8283: 	add	%r1, %r0, %r6
"10000100000001001101100000000000",	-- 8284: 	add	%r27, %r0, %r4
"00111111111111100000000000000101",	-- 8285: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 8286: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 8287: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 8288: 	jalr	%r26
"10101011110111100000000000000110",	-- 8289: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 8290: 	lw	%ra, [%sp + 5]
	-- bneq_cont.9215:
"11001100000000010000000000000001",	-- 8291: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 8292: 	lw	%r2, [%sp + 4]
"00101000010000010000000000000010",	-- 8293: 	bneq	%r2, %r1, bneq_else.9216
"01010100000000000010000001110110",	-- 8294: 	j	bneq_cont.9217
	-- bneq_else.9216:
"11001100000000010000000000000001",	-- 8295: 	lli	%r1, 1
"00111011110000110000000000000011",	-- 8296: 	lw	%r3, [%sp + 3]
"10000100011000010000100000000000",	-- 8297: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 8298: 	lw	%r1, [%r1 + 0]
"00111011110001000000000000000001",	-- 8299: 	lw	%r4, [%sp + 1]
"00111011110001010000000000000000",	-- 8300: 	lw	%r5, [%sp + 0]
"00111011110110110000000000000010",	-- 8301: 	lw	%r27, [%sp + 2]
"10000100000001010001100000000000",	-- 8302: 	add	%r3, %r0, %r5
"10000100000001000001000000000000",	-- 8303: 	add	%r2, %r0, %r4
"00111111111111100000000000000101",	-- 8304: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 8305: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 8306: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 8307: 	jalr	%r26
"10101011110111100000000000000110",	-- 8308: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 8309: 	lw	%ra, [%sp + 5]
	-- bneq_cont.9217:
"11001100000000010000000000000010",	-- 8310: 	lli	%r1, 2
"00111011110000100000000000000100",	-- 8311: 	lw	%r2, [%sp + 4]
"00101000010000010000000000000010",	-- 8312: 	bneq	%r2, %r1, bneq_else.9218
"01010100000000000010000010001001",	-- 8313: 	j	bneq_cont.9219
	-- bneq_else.9218:
"11001100000000010000000000000010",	-- 8314: 	lli	%r1, 2
"00111011110000110000000000000011",	-- 8315: 	lw	%r3, [%sp + 3]
"10000100011000010000100000000000",	-- 8316: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 8317: 	lw	%r1, [%r1 + 0]
"00111011110001000000000000000001",	-- 8318: 	lw	%r4, [%sp + 1]
"00111011110001010000000000000000",	-- 8319: 	lw	%r5, [%sp + 0]
"00111011110110110000000000000010",	-- 8320: 	lw	%r27, [%sp + 2]
"10000100000001010001100000000000",	-- 8321: 	add	%r3, %r0, %r5
"10000100000001000001000000000000",	-- 8322: 	add	%r2, %r0, %r4
"00111111111111100000000000000101",	-- 8323: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 8324: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 8325: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 8326: 	jalr	%r26
"10101011110111100000000000000110",	-- 8327: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 8328: 	lw	%ra, [%sp + 5]
	-- bneq_cont.9219:
"11001100000000010000000000000011",	-- 8329: 	lli	%r1, 3
"00111011110000100000000000000100",	-- 8330: 	lw	%r2, [%sp + 4]
"00101000010000010000000000000010",	-- 8331: 	bneq	%r2, %r1, bneq_else.9220
"01010100000000000010000010011100",	-- 8332: 	j	bneq_cont.9221
	-- bneq_else.9220:
"11001100000000010000000000000011",	-- 8333: 	lli	%r1, 3
"00111011110000110000000000000011",	-- 8334: 	lw	%r3, [%sp + 3]
"10000100011000010000100000000000",	-- 8335: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 8336: 	lw	%r1, [%r1 + 0]
"00111011110001000000000000000001",	-- 8337: 	lw	%r4, [%sp + 1]
"00111011110001010000000000000000",	-- 8338: 	lw	%r5, [%sp + 0]
"00111011110110110000000000000010",	-- 8339: 	lw	%r27, [%sp + 2]
"10000100000001010001100000000000",	-- 8340: 	add	%r3, %r0, %r5
"10000100000001000001000000000000",	-- 8341: 	add	%r2, %r0, %r4
"00111111111111100000000000000101",	-- 8342: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 8343: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 8344: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 8345: 	jalr	%r26
"10101011110111100000000000000110",	-- 8346: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 8347: 	lw	%ra, [%sp + 5]
	-- bneq_cont.9221:
"11001100000000010000000000000100",	-- 8348: 	lli	%r1, 4
"00111011110000100000000000000100",	-- 8349: 	lw	%r2, [%sp + 4]
"00101000010000010000000000000010",	-- 8350: 	bneq	%r2, %r1, bneq_else.9222
"01001111111000000000000000000000",	-- 8351: 	jr	%ra
	-- bneq_else.9222:
"11001100000000010000000000000100",	-- 8352: 	lli	%r1, 4
"00111011110000100000000000000011",	-- 8353: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 8354: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8355: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000000001",	-- 8356: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 8357: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000010",	-- 8358: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 8359: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8360: 	jr	%r26
	-- calc_diffuse_using_1point.2925:
"00111011011000110000000000000011",	-- 8361: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 8362: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 8363: 	lw	%r5, [%r27 + 1]
"00111100100111100000000000000000",	-- 8364: 	sw	%r4, [%sp + 0]
"00111100011111100000000000000001",	-- 8365: 	sw	%r3, [%sp + 1]
"00111100101111100000000000000010",	-- 8366: 	sw	%r5, [%sp + 2]
"00111100010111100000000000000011",	-- 8367: 	sw	%r2, [%sp + 3]
"00111100001111100000000000000100",	-- 8368: 	sw	%r1, [%sp + 4]
"00111111111111100000000000000101",	-- 8369: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 8370: 	addi	%sp, %sp, 6
"01011000000000000000011010101100",	-- 8371: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000000110",	-- 8372: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 8373: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000100",	-- 8374: 	lw	%r2, [%sp + 4]
"00111100001111100000000000000101",	-- 8375: 	sw	%r1, [%sp + 5]
"10000100000000100000100000000000",	-- 8376: 	add	%r1, %r0, %r2
"00111111111111100000000000000110",	-- 8377: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8378: 	addi	%sp, %sp, 7
"01011000000000000000011010111000",	-- 8379: 	jal	p_nvectors.2681
"10101011110111100000000000000111",	-- 8380: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8381: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000100",	-- 8382: 	lw	%r2, [%sp + 4]
"00111100001111100000000000000110",	-- 8383: 	sw	%r1, [%sp + 6]
"10000100000000100000100000000000",	-- 8384: 	add	%r1, %r0, %r2
"00111111111111100000000000000111",	-- 8385: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 8386: 	addi	%sp, %sp, 8
"01011000000000000000011010100100",	-- 8387: 	jal	p_intersection_points.2666
"10101011110111100000000000001000",	-- 8388: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8389: 	lw	%ra, [%sp + 7]
"00111011110000100000000000000100",	-- 8390: 	lw	%r2, [%sp + 4]
"00111100001111100000000000000111",	-- 8391: 	sw	%r1, [%sp + 7]
"10000100000000100000100000000000",	-- 8392: 	add	%r1, %r0, %r2
"00111111111111100000000000001000",	-- 8393: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 8394: 	addi	%sp, %sp, 9
"01011000000000000000011010101010",	-- 8395: 	jal	p_energy.2672
"10101011110111100000000000001001",	-- 8396: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 8397: 	lw	%ra, [%sp + 8]
"00111011110000100000000000000011",	-- 8398: 	lw	%r2, [%sp + 3]
"00111011110000110000000000000101",	-- 8399: 	lw	%r3, [%sp + 5]
"10000100011000100001100000000000",	-- 8400: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 8401: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000000010",	-- 8402: 	lw	%r4, [%sp + 2]
"00111100001111100000000000001000",	-- 8403: 	sw	%r1, [%sp + 8]
"10000100000000110001000000000000",	-- 8404: 	add	%r2, %r0, %r3
"10000100000001000000100000000000",	-- 8405: 	add	%r1, %r0, %r4
"00111111111111100000000000001001",	-- 8406: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 8407: 	addi	%sp, %sp, 10
"01011000000000000000010100111011",	-- 8408: 	jal	veccpy.2586
"10101011110111100000000000001010",	-- 8409: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 8410: 	lw	%ra, [%sp + 9]
"00111011110000010000000000000100",	-- 8411: 	lw	%r1, [%sp + 4]
"00111111111111100000000000001001",	-- 8412: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 8413: 	addi	%sp, %sp, 10
"01011000000000000000011010101110",	-- 8414: 	jal	p_group_id.2676
"10101011110111100000000000001010",	-- 8415: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 8416: 	lw	%ra, [%sp + 9]
"00111011110000100000000000000011",	-- 8417: 	lw	%r2, [%sp + 3]
"00111011110000110000000000000110",	-- 8418: 	lw	%r3, [%sp + 6]
"10000100011000100001100000000000",	-- 8419: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 8420: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000000111",	-- 8421: 	lw	%r4, [%sp + 7]
"10000100100000100010000000000000",	-- 8422: 	add	%r4, %r4, %r2
"00111000100001000000000000000000",	-- 8423: 	lw	%r4, [%r4 + 0]
"00111011110110110000000000000001",	-- 8424: 	lw	%r27, [%sp + 1]
"10000100000000110001000000000000",	-- 8425: 	add	%r2, %r0, %r3
"10000100000001000001100000000000",	-- 8426: 	add	%r3, %r0, %r4
"00111111111111100000000000001001",	-- 8427: 	sw	%ra, [%sp + 9]
"00111011011110100000000000000000",	-- 8428: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001010",	-- 8429: 	addi	%sp, %sp, 10
"01010011010000000000000000000000",	-- 8430: 	jalr	%r26
"10101011110111100000000000001010",	-- 8431: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 8432: 	lw	%ra, [%sp + 9]
"00111011110000010000000000000011",	-- 8433: 	lw	%r1, [%sp + 3]
"00111011110000100000000000001000",	-- 8434: 	lw	%r2, [%sp + 8]
"10000100010000010000100000000000",	-- 8435: 	add	%r1, %r2, %r1
"00111000001000100000000000000000",	-- 8436: 	lw	%r2, [%r1 + 0]
"00111011110000010000000000000000",	-- 8437: 	lw	%r1, [%sp + 0]
"00111011110000110000000000000010",	-- 8438: 	lw	%r3, [%sp + 2]
"01010100000000000000011000100011",	-- 8439: 	j	vecaccumv.2618
	-- calc_diffuse_using_5points.2928:
"00111011011001100000000000000010",	-- 8440: 	lw	%r6, [%r27 + 2]
"00111011011001110000000000000001",	-- 8441: 	lw	%r7, [%r27 + 1]
"10000100010000010001000000000000",	-- 8442: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 8443: 	lw	%r2, [%r2 + 0]
"00111100110111100000000000000000",	-- 8444: 	sw	%r6, [%sp + 0]
"00111100111111100000000000000001",	-- 8445: 	sw	%r7, [%sp + 1]
"00111100101111100000000000000010",	-- 8446: 	sw	%r5, [%sp + 2]
"00111100100111100000000000000011",	-- 8447: 	sw	%r4, [%sp + 3]
"00111100011111100000000000000100",	-- 8448: 	sw	%r3, [%sp + 4]
"00111100001111100000000000000101",	-- 8449: 	sw	%r1, [%sp + 5]
"10000100000000100000100000000000",	-- 8450: 	add	%r1, %r0, %r2
"00111111111111100000000000000110",	-- 8451: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8452: 	addi	%sp, %sp, 7
"01011000000000000000011010101100",	-- 8453: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000000111",	-- 8454: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8455: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000001",	-- 8456: 	lli	%r2, 1
"00111011110000110000000000000101",	-- 8457: 	lw	%r3, [%sp + 5]
"10001000011000100001000000000000",	-- 8458: 	sub	%r2, %r3, %r2
"00111011110001000000000000000100",	-- 8459: 	lw	%r4, [%sp + 4]
"10000100100000100001000000000000",	-- 8460: 	add	%r2, %r4, %r2
"00111000010000100000000000000000",	-- 8461: 	lw	%r2, [%r2 + 0]
"00111100001111100000000000000110",	-- 8462: 	sw	%r1, [%sp + 6]
"10000100000000100000100000000000",	-- 8463: 	add	%r1, %r0, %r2
"00111111111111100000000000000111",	-- 8464: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 8465: 	addi	%sp, %sp, 8
"01011000000000000000011010101100",	-- 8466: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000001000",	-- 8467: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8468: 	lw	%ra, [%sp + 7]
"00111011110000100000000000000101",	-- 8469: 	lw	%r2, [%sp + 5]
"00111011110000110000000000000100",	-- 8470: 	lw	%r3, [%sp + 4]
"10000100011000100010000000000000",	-- 8471: 	add	%r4, %r3, %r2
"00111000100001000000000000000000",	-- 8472: 	lw	%r4, [%r4 + 0]
"00111100001111100000000000000111",	-- 8473: 	sw	%r1, [%sp + 7]
"10000100000001000000100000000000",	-- 8474: 	add	%r1, %r0, %r4
"00111111111111100000000000001000",	-- 8475: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 8476: 	addi	%sp, %sp, 9
"01011000000000000000011010101100",	-- 8477: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000001001",	-- 8478: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 8479: 	lw	%ra, [%sp + 8]
"11001100000000100000000000000001",	-- 8480: 	lli	%r2, 1
"00111011110000110000000000000101",	-- 8481: 	lw	%r3, [%sp + 5]
"10000100011000100001000000000000",	-- 8482: 	add	%r2, %r3, %r2
"00111011110001000000000000000100",	-- 8483: 	lw	%r4, [%sp + 4]
"10000100100000100001000000000000",	-- 8484: 	add	%r2, %r4, %r2
"00111000010000100000000000000000",	-- 8485: 	lw	%r2, [%r2 + 0]
"00111100001111100000000000001000",	-- 8486: 	sw	%r1, [%sp + 8]
"10000100000000100000100000000000",	-- 8487: 	add	%r1, %r0, %r2
"00111111111111100000000000001001",	-- 8488: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 8489: 	addi	%sp, %sp, 10
"01011000000000000000011010101100",	-- 8490: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000001010",	-- 8491: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 8492: 	lw	%ra, [%sp + 9]
"00111011110000100000000000000101",	-- 8493: 	lw	%r2, [%sp + 5]
"00111011110000110000000000000011",	-- 8494: 	lw	%r3, [%sp + 3]
"10000100011000100001100000000000",	-- 8495: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 8496: 	lw	%r3, [%r3 + 0]
"00111100001111100000000000001001",	-- 8497: 	sw	%r1, [%sp + 9]
"10000100000000110000100000000000",	-- 8498: 	add	%r1, %r0, %r3
"00111111111111100000000000001010",	-- 8499: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 8500: 	addi	%sp, %sp, 11
"01011000000000000000011010101100",	-- 8501: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000001011",	-- 8502: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 8503: 	lw	%ra, [%sp + 10]
"00111011110000100000000000000010",	-- 8504: 	lw	%r2, [%sp + 2]
"00111011110000110000000000000110",	-- 8505: 	lw	%r3, [%sp + 6]
"10000100011000100001100000000000",	-- 8506: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 8507: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000000001",	-- 8508: 	lw	%r4, [%sp + 1]
"00111100001111100000000000001010",	-- 8509: 	sw	%r1, [%sp + 10]
"10000100000000110001000000000000",	-- 8510: 	add	%r2, %r0, %r3
"10000100000001000000100000000000",	-- 8511: 	add	%r1, %r0, %r4
"00111111111111100000000000001011",	-- 8512: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8513: 	addi	%sp, %sp, 12
"01011000000000000000010100111011",	-- 8514: 	jal	veccpy.2586
"10101011110111100000000000001100",	-- 8515: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8516: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000010",	-- 8517: 	lw	%r1, [%sp + 2]
"00111011110000100000000000000111",	-- 8518: 	lw	%r2, [%sp + 7]
"10000100010000010001000000000000",	-- 8519: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 8520: 	lw	%r2, [%r2 + 0]
"00111011110000110000000000000001",	-- 8521: 	lw	%r3, [%sp + 1]
"10000100000000110000100000000000",	-- 8522: 	add	%r1, %r0, %r3
"00111111111111100000000000001011",	-- 8523: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8524: 	addi	%sp, %sp, 12
"01011000000000000000010111101110",	-- 8525: 	jal	vecadd.2609
"10101011110111100000000000001100",	-- 8526: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8527: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000010",	-- 8528: 	lw	%r1, [%sp + 2]
"00111011110000100000000000001000",	-- 8529: 	lw	%r2, [%sp + 8]
"10000100010000010001000000000000",	-- 8530: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 8531: 	lw	%r2, [%r2 + 0]
"00111011110000110000000000000001",	-- 8532: 	lw	%r3, [%sp + 1]
"10000100000000110000100000000000",	-- 8533: 	add	%r1, %r0, %r3
"00111111111111100000000000001011",	-- 8534: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8535: 	addi	%sp, %sp, 12
"01011000000000000000010111101110",	-- 8536: 	jal	vecadd.2609
"10101011110111100000000000001100",	-- 8537: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8538: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000010",	-- 8539: 	lw	%r1, [%sp + 2]
"00111011110000100000000000001001",	-- 8540: 	lw	%r2, [%sp + 9]
"10000100010000010001000000000000",	-- 8541: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 8542: 	lw	%r2, [%r2 + 0]
"00111011110000110000000000000001",	-- 8543: 	lw	%r3, [%sp + 1]
"10000100000000110000100000000000",	-- 8544: 	add	%r1, %r0, %r3
"00111111111111100000000000001011",	-- 8545: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8546: 	addi	%sp, %sp, 12
"01011000000000000000010111101110",	-- 8547: 	jal	vecadd.2609
"10101011110111100000000000001100",	-- 8548: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8549: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000010",	-- 8550: 	lw	%r1, [%sp + 2]
"00111011110000100000000000001010",	-- 8551: 	lw	%r2, [%sp + 10]
"10000100010000010001000000000000",	-- 8552: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 8553: 	lw	%r2, [%r2 + 0]
"00111011110000110000000000000001",	-- 8554: 	lw	%r3, [%sp + 1]
"10000100000000110000100000000000",	-- 8555: 	add	%r1, %r0, %r3
"00111111111111100000000000001011",	-- 8556: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8557: 	addi	%sp, %sp, 12
"01011000000000000000010111101110",	-- 8558: 	jal	vecadd.2609
"10101011110111100000000000001100",	-- 8559: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8560: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000101",	-- 8561: 	lw	%r1, [%sp + 5]
"00111011110000100000000000000100",	-- 8562: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 8563: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8564: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001011",	-- 8565: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8566: 	addi	%sp, %sp, 12
"01011000000000000000011010101010",	-- 8567: 	jal	p_energy.2672
"10101011110111100000000000001100",	-- 8568: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8569: 	lw	%ra, [%sp + 11]
"00111011110000100000000000000010",	-- 8570: 	lw	%r2, [%sp + 2]
"10000100001000100000100000000000",	-- 8571: 	add	%r1, %r1, %r2
"00111000001000100000000000000000",	-- 8572: 	lw	%r2, [%r1 + 0]
"00111011110000010000000000000000",	-- 8573: 	lw	%r1, [%sp + 0]
"00111011110000110000000000000001",	-- 8574: 	lw	%r3, [%sp + 1]
"01010100000000000000011000100011",	-- 8575: 	j	vecaccumv.2618
	-- do_without_neighbors.2934:
"00111011011000110000000000000001",	-- 8576: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000100",	-- 8577: 	lli	%r4, 4
"00110000010001000000000000101011",	-- 8578: 	bgt	%r2, %r4, bgt_else.9224
"00111111011111100000000000000000",	-- 8579: 	sw	%r27, [%sp + 0]
"00111100011111100000000000000001",	-- 8580: 	sw	%r3, [%sp + 1]
"00111100001111100000000000000010",	-- 8581: 	sw	%r1, [%sp + 2]
"00111100010111100000000000000011",	-- 8582: 	sw	%r2, [%sp + 3]
"00111111111111100000000000000100",	-- 8583: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 8584: 	addi	%sp, %sp, 5
"01011000000000000000011010100110",	-- 8585: 	jal	p_surface_ids.2668
"10101011110111100000000000000101",	-- 8586: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 8587: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000000",	-- 8588: 	lli	%r2, 0
"00111011110000110000000000000011",	-- 8589: 	lw	%r3, [%sp + 3]
"10000100001000110000100000000000",	-- 8590: 	add	%r1, %r1, %r3
"00111000001000010000000000000000",	-- 8591: 	lw	%r1, [%r1 + 0]
"00110000010000010000000000011100",	-- 8592: 	bgt	%r2, %r1, bgt_else.9225
"00111011110000010000000000000010",	-- 8593: 	lw	%r1, [%sp + 2]
"00111111111111100000000000000100",	-- 8594: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 8595: 	addi	%sp, %sp, 5
"01011000000000000000011010101000",	-- 8596: 	jal	p_calc_diffuse.2670
"10101011110111100000000000000101",	-- 8597: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 8598: 	lw	%ra, [%sp + 4]
"00111011110000100000000000000011",	-- 8599: 	lw	%r2, [%sp + 3]
"10000100001000100000100000000000",	-- 8600: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 8601: 	lw	%r1, [%r1 + 0]
"11001100000000110000000000000000",	-- 8602: 	lli	%r3, 0
"00101000001000110000000000000010",	-- 8603: 	bneq	%r1, %r3, bneq_else.9226
"01010100000000000010000110100101",	-- 8604: 	j	bneq_cont.9227
	-- bneq_else.9226:
"00111011110000010000000000000010",	-- 8605: 	lw	%r1, [%sp + 2]
"00111011110110110000000000000001",	-- 8606: 	lw	%r27, [%sp + 1]
"00111111111111100000000000000100",	-- 8607: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 8608: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 8609: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 8610: 	jalr	%r26
"10101011110111100000000000000101",	-- 8611: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 8612: 	lw	%ra, [%sp + 4]
	-- bneq_cont.9227:
"11001100000000010000000000000001",	-- 8613: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 8614: 	lw	%r2, [%sp + 3]
"10000100010000010001000000000000",	-- 8615: 	add	%r2, %r2, %r1
"00111011110000010000000000000010",	-- 8616: 	lw	%r1, [%sp + 2]
"00111011110110110000000000000000",	-- 8617: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 8618: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8619: 	jr	%r26
	-- bgt_else.9225:
"01001111111000000000000000000000",	-- 8620: 	jr	%ra
	-- bgt_else.9224:
"01001111111000000000000000000000",	-- 8621: 	jr	%ra
	-- neighbors_exist.2937:
"00111011011000110000000000000001",	-- 8622: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000001",	-- 8623: 	lli	%r4, 1
"10000100011001000010000000000000",	-- 8624: 	add	%r4, %r3, %r4
"00111000100001000000000000000000",	-- 8625: 	lw	%r4, [%r4 + 0]
"11001100000001010000000000000001",	-- 8626: 	lli	%r5, 1
"10000100010001010010100000000000",	-- 8627: 	add	%r5, %r2, %r5
"00110000100001010000000000000011",	-- 8628: 	bgt	%r4, %r5, bgt_else.9230
"11001100000000010000000000000000",	-- 8629: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8630: 	jr	%ra
	-- bgt_else.9230:
"11001100000001000000000000000000",	-- 8631: 	lli	%r4, 0
"00110000010001000000000000000011",	-- 8632: 	bgt	%r2, %r4, bgt_else.9231
"11001100000000010000000000000000",	-- 8633: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8634: 	jr	%ra
	-- bgt_else.9231:
"11001100000000100000000000000000",	-- 8635: 	lli	%r2, 0
"10000100011000100001000000000000",	-- 8636: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 8637: 	lw	%r2, [%r2 + 0]
"11001100000000110000000000000001",	-- 8638: 	lli	%r3, 1
"10000100001000110001100000000000",	-- 8639: 	add	%r3, %r1, %r3
"00110000010000110000000000000011",	-- 8640: 	bgt	%r2, %r3, bgt_else.9232
"11001100000000010000000000000000",	-- 8641: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8642: 	jr	%ra
	-- bgt_else.9232:
"11001100000000100000000000000000",	-- 8643: 	lli	%r2, 0
"00110000001000100000000000000011",	-- 8644: 	bgt	%r1, %r2, bgt_else.9233
"11001100000000010000000000000000",	-- 8645: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8646: 	jr	%ra
	-- bgt_else.9233:
"11001100000000010000000000000001",	-- 8647: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 8648: 	jr	%ra
	-- get_surface_id.2941:
"00111100010111100000000000000000",	-- 8649: 	sw	%r2, [%sp + 0]
"00111111111111100000000000000001",	-- 8650: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8651: 	addi	%sp, %sp, 2
"01011000000000000000011010100110",	-- 8652: 	jal	p_surface_ids.2668
"10101011110111100000000000000010",	-- 8653: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8654: 	lw	%ra, [%sp + 1]
"00111011110000100000000000000000",	-- 8655: 	lw	%r2, [%sp + 0]
"10000100001000100000100000000000",	-- 8656: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 8657: 	lw	%r1, [%r1 + 0]
"01001111111000000000000000000000",	-- 8658: 	jr	%ra
	-- neighbors_are_available.2944:
"10000100011000010011000000000000",	-- 8659: 	add	%r6, %r3, %r1
"00111000110001100000000000000000",	-- 8660: 	lw	%r6, [%r6 + 0]
"00111100011111100000000000000000",	-- 8661: 	sw	%r3, [%sp + 0]
"00111100100111100000000000000001",	-- 8662: 	sw	%r4, [%sp + 1]
"00111100101111100000000000000010",	-- 8663: 	sw	%r5, [%sp + 2]
"00111100001111100000000000000011",	-- 8664: 	sw	%r1, [%sp + 3]
"00111100010111100000000000000100",	-- 8665: 	sw	%r2, [%sp + 4]
"10000100000001010001000000000000",	-- 8666: 	add	%r2, %r0, %r5
"10000100000001100000100000000000",	-- 8667: 	add	%r1, %r0, %r6
"00111111111111100000000000000101",	-- 8668: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 8669: 	addi	%sp, %sp, 6
"01011000000000000010000111001001",	-- 8670: 	jal	get_surface_id.2941
"10101011110111100000000000000110",	-- 8671: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 8672: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000011",	-- 8673: 	lw	%r2, [%sp + 3]
"00111011110000110000000000000100",	-- 8674: 	lw	%r3, [%sp + 4]
"10000100011000100001100000000000",	-- 8675: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 8676: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000000010",	-- 8677: 	lw	%r4, [%sp + 2]
"00111100001111100000000000000101",	-- 8678: 	sw	%r1, [%sp + 5]
"10000100000001000001000000000000",	-- 8679: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 8680: 	add	%r1, %r0, %r3
"00111111111111100000000000000110",	-- 8681: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8682: 	addi	%sp, %sp, 7
"01011000000000000010000111001001",	-- 8683: 	jal	get_surface_id.2941
"10101011110111100000000000000111",	-- 8684: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8685: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000101",	-- 8686: 	lw	%r2, [%sp + 5]
"00101000001000100000000000110101",	-- 8687: 	bneq	%r1, %r2, bneq_else.9234
"00111011110000010000000000000011",	-- 8688: 	lw	%r1, [%sp + 3]
"00111011110000110000000000000001",	-- 8689: 	lw	%r3, [%sp + 1]
"10000100011000010001100000000000",	-- 8690: 	add	%r3, %r3, %r1
"00111000011000110000000000000000",	-- 8691: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000000010",	-- 8692: 	lw	%r4, [%sp + 2]
"10000100000001000001000000000000",	-- 8693: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 8694: 	add	%r1, %r0, %r3
"00111111111111100000000000000110",	-- 8695: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8696: 	addi	%sp, %sp, 7
"01011000000000000010000111001001",	-- 8697: 	jal	get_surface_id.2941
"10101011110111100000000000000111",	-- 8698: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8699: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000101",	-- 8700: 	lw	%r2, [%sp + 5]
"00101000001000100000000000100101",	-- 8701: 	bneq	%r1, %r2, bneq_else.9235
"11001100000000010000000000000001",	-- 8702: 	lli	%r1, 1
"00111011110000110000000000000011",	-- 8703: 	lw	%r3, [%sp + 3]
"10001000011000010000100000000000",	-- 8704: 	sub	%r1, %r3, %r1
"00111011110001000000000000000000",	-- 8705: 	lw	%r4, [%sp + 0]
"10000100100000010000100000000000",	-- 8706: 	add	%r1, %r4, %r1
"00111000001000010000000000000000",	-- 8707: 	lw	%r1, [%r1 + 0]
"00111011110001010000000000000010",	-- 8708: 	lw	%r5, [%sp + 2]
"10000100000001010001000000000000",	-- 8709: 	add	%r2, %r0, %r5
"00111111111111100000000000000110",	-- 8710: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8711: 	addi	%sp, %sp, 7
"01011000000000000010000111001001",	-- 8712: 	jal	get_surface_id.2941
"10101011110111100000000000000111",	-- 8713: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8714: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000101",	-- 8715: 	lw	%r2, [%sp + 5]
"00101000001000100000000000010100",	-- 8716: 	bneq	%r1, %r2, bneq_else.9236
"11001100000000010000000000000001",	-- 8717: 	lli	%r1, 1
"00111011110000110000000000000011",	-- 8718: 	lw	%r3, [%sp + 3]
"10000100011000010000100000000000",	-- 8719: 	add	%r1, %r3, %r1
"00111011110000110000000000000000",	-- 8720: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 8721: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 8722: 	lw	%r1, [%r1 + 0]
"00111011110000110000000000000010",	-- 8723: 	lw	%r3, [%sp + 2]
"10000100000000110001000000000000",	-- 8724: 	add	%r2, %r0, %r3
"00111111111111100000000000000110",	-- 8725: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8726: 	addi	%sp, %sp, 7
"01011000000000000010000111001001",	-- 8727: 	jal	get_surface_id.2941
"10101011110111100000000000000111",	-- 8728: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8729: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000101",	-- 8730: 	lw	%r2, [%sp + 5]
"00101000001000100000000000000011",	-- 8731: 	bneq	%r1, %r2, bneq_else.9237
"11001100000000010000000000000001",	-- 8732: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 8733: 	jr	%ra
	-- bneq_else.9237:
"11001100000000010000000000000000",	-- 8734: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8735: 	jr	%ra
	-- bneq_else.9236:
"11001100000000010000000000000000",	-- 8736: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8737: 	jr	%ra
	-- bneq_else.9235:
"11001100000000010000000000000000",	-- 8738: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8739: 	jr	%ra
	-- bneq_else.9234:
"11001100000000010000000000000000",	-- 8740: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8741: 	jr	%ra
	-- try_exploit_neighbors.2950:
"00111011011001110000000000000010",	-- 8742: 	lw	%r7, [%r27 + 2]
"00111011011010000000000000000001",	-- 8743: 	lw	%r8, [%r27 + 1]
"10000100100000010100100000000000",	-- 8744: 	add	%r9, %r4, %r1
"00111001001010010000000000000000",	-- 8745: 	lw	%r9, [%r9 + 0]
"11001100000010100000000000000100",	-- 8746: 	lli	%r10, 4
"00110000110010100000000001001101",	-- 8747: 	bgt	%r6, %r10, bgt_else.9238
"11001100000010100000000000000000",	-- 8748: 	lli	%r10, 0
"00111100010111100000000000000000",	-- 8749: 	sw	%r2, [%sp + 0]
"00111111011111100000000000000001",	-- 8750: 	sw	%r27, [%sp + 1]
"00111101000111100000000000000010",	-- 8751: 	sw	%r8, [%sp + 2]
"00111101001111100000000000000011",	-- 8752: 	sw	%r9, [%sp + 3]
"00111100111111100000000000000100",	-- 8753: 	sw	%r7, [%sp + 4]
"00111100110111100000000000000101",	-- 8754: 	sw	%r6, [%sp + 5]
"00111100101111100000000000000110",	-- 8755: 	sw	%r5, [%sp + 6]
"00111100100111100000000000000111",	-- 8756: 	sw	%r4, [%sp + 7]
"00111100011111100000000000001000",	-- 8757: 	sw	%r3, [%sp + 8]
"00111100001111100000000000001001",	-- 8758: 	sw	%r1, [%sp + 9]
"00111101010111100000000000001010",	-- 8759: 	sw	%r10, [%sp + 10]
"10000100000001100001000000000000",	-- 8760: 	add	%r2, %r0, %r6
"10000100000010010000100000000000",	-- 8761: 	add	%r1, %r0, %r9
"00111111111111100000000000001011",	-- 8762: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8763: 	addi	%sp, %sp, 12
"01011000000000000010000111001001",	-- 8764: 	jal	get_surface_id.2941
"10101011110111100000000000001100",	-- 8765: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8766: 	lw	%ra, [%sp + 11]
"00111011110000100000000000001010",	-- 8767: 	lw	%r2, [%sp + 10]
"00110000010000010000000000110111",	-- 8768: 	bgt	%r2, %r1, bgt_else.9239
"00111011110000010000000000001001",	-- 8769: 	lw	%r1, [%sp + 9]
"00111011110000100000000000001000",	-- 8770: 	lw	%r2, [%sp + 8]
"00111011110000110000000000000111",	-- 8771: 	lw	%r3, [%sp + 7]
"00111011110001000000000000000110",	-- 8772: 	lw	%r4, [%sp + 6]
"00111011110001010000000000000101",	-- 8773: 	lw	%r5, [%sp + 5]
"00111111111111100000000000001011",	-- 8774: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8775: 	addi	%sp, %sp, 12
"01011000000000000010000111010011",	-- 8776: 	jal	neighbors_are_available.2944
"10101011110111100000000000001100",	-- 8777: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8778: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 8779: 	lli	%r2, 0
"00101000001000100000000000001001",	-- 8780: 	bneq	%r1, %r2, bneq_else.9240
"00111011110000010000000000001001",	-- 8781: 	lw	%r1, [%sp + 9]
"00111011110000100000000000000111",	-- 8782: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 8783: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8784: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000000101",	-- 8785: 	lw	%r2, [%sp + 5]
"00111011110110110000000000000100",	-- 8786: 	lw	%r27, [%sp + 4]
"00111011011110100000000000000000",	-- 8787: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8788: 	jr	%r26
	-- bneq_else.9240:
"00111011110000010000000000000011",	-- 8789: 	lw	%r1, [%sp + 3]
"00111111111111100000000000001011",	-- 8790: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8791: 	addi	%sp, %sp, 12
"01011000000000000000011010101000",	-- 8792: 	jal	p_calc_diffuse.2670
"10101011110111100000000000001100",	-- 8793: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8794: 	lw	%ra, [%sp + 11]
"00111011110001010000000000000101",	-- 8795: 	lw	%r5, [%sp + 5]
"10000100001001010000100000000000",	-- 8796: 	add	%r1, %r1, %r5
"00111000001000010000000000000000",	-- 8797: 	lw	%r1, [%r1 + 0]
"11001100000000100000000000000000",	-- 8798: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 8799: 	bneq	%r1, %r2, bneq_else.9241
"01010100000000000010001001101100",	-- 8800: 	j	bneq_cont.9242
	-- bneq_else.9241:
"00111011110000010000000000001001",	-- 8801: 	lw	%r1, [%sp + 9]
"00111011110000100000000000001000",	-- 8802: 	lw	%r2, [%sp + 8]
"00111011110000110000000000000111",	-- 8803: 	lw	%r3, [%sp + 7]
"00111011110001000000000000000110",	-- 8804: 	lw	%r4, [%sp + 6]
"00111011110110110000000000000010",	-- 8805: 	lw	%r27, [%sp + 2]
"00111111111111100000000000001011",	-- 8806: 	sw	%ra, [%sp + 11]
"00111011011110100000000000000000",	-- 8807: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001100",	-- 8808: 	addi	%sp, %sp, 12
"01010011010000000000000000000000",	-- 8809: 	jalr	%r26
"10101011110111100000000000001100",	-- 8810: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8811: 	lw	%ra, [%sp + 11]
	-- bneq_cont.9242:
"11001100000000010000000000000001",	-- 8812: 	lli	%r1, 1
"00111011110000100000000000000101",	-- 8813: 	lw	%r2, [%sp + 5]
"10000100010000010011000000000000",	-- 8814: 	add	%r6, %r2, %r1
"00111011110000010000000000001001",	-- 8815: 	lw	%r1, [%sp + 9]
"00111011110000100000000000000000",	-- 8816: 	lw	%r2, [%sp + 0]
"00111011110000110000000000001000",	-- 8817: 	lw	%r3, [%sp + 8]
"00111011110001000000000000000111",	-- 8818: 	lw	%r4, [%sp + 7]
"00111011110001010000000000000110",	-- 8819: 	lw	%r5, [%sp + 6]
"00111011110110110000000000000001",	-- 8820: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 8821: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8822: 	jr	%r26
	-- bgt_else.9239:
"01001111111000000000000000000000",	-- 8823: 	jr	%ra
	-- bgt_else.9238:
"01001111111000000000000000000000",	-- 8824: 	jr	%ra
	-- write_ppm_header.2957:
"00111011011000010000000000000001",	-- 8825: 	lw	%r1, [%r27 + 1]
"11001100000000100000000001010000",	-- 8826: 	lli	%r2, 80
"00111100001111100000000000000000",	-- 8827: 	sw	%r1, [%sp + 0]
"10000100000000100000100000000000",	-- 8828: 	add	%r1, %r0, %r2
"00111111111111100000000000000001",	-- 8829: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8830: 	addi	%sp, %sp, 2
"01011000000000000010101000011000",	-- 8831: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8832: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8833: 	lw	%ra, [%sp + 1]
"11001100000000010000000000110011",	-- 8834: 	lli	%r1, 51
"00111111111111100000000000000001",	-- 8835: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8836: 	addi	%sp, %sp, 2
"01011000000000000010101000011000",	-- 8837: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8838: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8839: 	lw	%ra, [%sp + 1]
"11001100000000010000000000001010",	-- 8840: 	lli	%r1, 10
"00111111111111100000000000000001",	-- 8841: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8842: 	addi	%sp, %sp, 2
"01011000000000000010101000011000",	-- 8843: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8844: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8845: 	lw	%ra, [%sp + 1]
"11001100000000010000000000000000",	-- 8846: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 8847: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 8848: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8849: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000000001",	-- 8850: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8851: 	addi	%sp, %sp, 2
"01011000000000000000010000000000",	-- 8852: 	jal	print_int.2514
"10101011110111100000000000000010",	-- 8853: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8854: 	lw	%ra, [%sp + 1]
"11001100000000010000000000100000",	-- 8855: 	lli	%r1, 32
"00111111111111100000000000000001",	-- 8856: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8857: 	addi	%sp, %sp, 2
"01011000000000000010101000011000",	-- 8858: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8859: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8860: 	lw	%ra, [%sp + 1]
"11001100000000010000000000000001",	-- 8861: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 8862: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 8863: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8864: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000000001",	-- 8865: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8866: 	addi	%sp, %sp, 2
"01011000000000000000010000000000",	-- 8867: 	jal	print_int.2514
"10101011110111100000000000000010",	-- 8868: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8869: 	lw	%ra, [%sp + 1]
"11001100000000010000000000100000",	-- 8870: 	lli	%r1, 32
"00111111111111100000000000000001",	-- 8871: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8872: 	addi	%sp, %sp, 2
"01011000000000000010101000011000",	-- 8873: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8874: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8875: 	lw	%ra, [%sp + 1]
"11001100000000010000000011111111",	-- 8876: 	lli	%r1, 255
"00111111111111100000000000000001",	-- 8877: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8878: 	addi	%sp, %sp, 2
"01011000000000000000010000000000",	-- 8879: 	jal	print_int.2514
"10101011110111100000000000000010",	-- 8880: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8881: 	lw	%ra, [%sp + 1]
"11001100000000010000000000001010",	-- 8882: 	lli	%r1, 10
"01010100000000000010101000011000",	-- 8883: 	j	yj_print_char
	-- write_rgb_element.2959:
"00111111111111100000000000000000",	-- 8884: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 8885: 	addi	%sp, %sp, 1
"01011000000000000010101000101100",	-- 8886: 	jal	yj_int_of_float
"10101011110111100000000000000001",	-- 8887: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 8888: 	lw	%ra, [%sp + 0]
"11001100000000100000000011111111",	-- 8889: 	lli	%r2, 255
"00110000001000100000000000000110",	-- 8890: 	bgt	%r1, %r2, bgt_else.9245
"11001100000000100000000000000000",	-- 8891: 	lli	%r2, 0
"00110000010000010000000000000010",	-- 8892: 	bgt	%r2, %r1, bgt_else.9247
"01010100000000000010001010111111",	-- 8893: 	j	bgt_cont.9248
	-- bgt_else.9247:
"11001100000000010000000000000000",	-- 8894: 	lli	%r1, 0
	-- bgt_cont.9248:
"01010100000000000010001011000001",	-- 8895: 	j	bgt_cont.9246
	-- bgt_else.9245:
"11001100000000010000000011111111",	-- 8896: 	lli	%r1, 255
	-- bgt_cont.9246:
"01010100000000000000010000000000",	-- 8897: 	j	print_int.2514
	-- write_rgb.2961:
"00111011011000010000000000000001",	-- 8898: 	lw	%r1, [%r27 + 1]
"11001100000000100000000000000000",	-- 8899: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 8900: 	add	%r2, %r1, %r2
"10010000010000000000000000000000",	-- 8901: 	lf	%f0, [%r2 + 0]
"00111100001111100000000000000000",	-- 8902: 	sw	%r1, [%sp + 0]
"00111111111111100000000000000001",	-- 8903: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8904: 	addi	%sp, %sp, 2
"01011000000000000010001010110100",	-- 8905: 	jal	write_rgb_element.2959
"10101011110111100000000000000010",	-- 8906: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8907: 	lw	%ra, [%sp + 1]
"11001100000000010000000000100000",	-- 8908: 	lli	%r1, 32
"00111111111111100000000000000001",	-- 8909: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8910: 	addi	%sp, %sp, 2
"01011000000000000010101000011000",	-- 8911: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8912: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8913: 	lw	%ra, [%sp + 1]
"11001100000000010000000000000001",	-- 8914: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 8915: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 8916: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 8917: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000000001",	-- 8918: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8919: 	addi	%sp, %sp, 2
"01011000000000000010001010110100",	-- 8920: 	jal	write_rgb_element.2959
"10101011110111100000000000000010",	-- 8921: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8922: 	lw	%ra, [%sp + 1]
"11001100000000010000000000100000",	-- 8923: 	lli	%r1, 32
"00111111111111100000000000000001",	-- 8924: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8925: 	addi	%sp, %sp, 2
"01011000000000000010101000011000",	-- 8926: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8927: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8928: 	lw	%ra, [%sp + 1]
"11001100000000010000000000000010",	-- 8929: 	lli	%r1, 2
"00111011110000100000000000000000",	-- 8930: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 8931: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 8932: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000000001",	-- 8933: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8934: 	addi	%sp, %sp, 2
"01011000000000000010001010110100",	-- 8935: 	jal	write_rgb_element.2959
"10101011110111100000000000000010",	-- 8936: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8937: 	lw	%ra, [%sp + 1]
"11001100000000010000000000001010",	-- 8938: 	lli	%r1, 10
"01010100000000000010101000011000",	-- 8939: 	j	yj_print_char
	-- pretrace_diffuse_rays.2963:
"00111011011000110000000000000011",	-- 8940: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 8941: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 8942: 	lw	%r5, [%r27 + 1]
"11001100000001100000000000000100",	-- 8943: 	lli	%r6, 4
"00110000010001100000000001100010",	-- 8944: 	bgt	%r2, %r6, bgt_else.9249
"00111111011111100000000000000000",	-- 8945: 	sw	%r27, [%sp + 0]
"00111100011111100000000000000001",	-- 8946: 	sw	%r3, [%sp + 1]
"00111100100111100000000000000010",	-- 8947: 	sw	%r4, [%sp + 2]
"00111100101111100000000000000011",	-- 8948: 	sw	%r5, [%sp + 3]
"00111100010111100000000000000100",	-- 8949: 	sw	%r2, [%sp + 4]
"00111100001111100000000000000101",	-- 8950: 	sw	%r1, [%sp + 5]
"00111111111111100000000000000110",	-- 8951: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8952: 	addi	%sp, %sp, 7
"01011000000000000010000111001001",	-- 8953: 	jal	get_surface_id.2941
"10101011110111100000000000000111",	-- 8954: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8955: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 8956: 	lli	%r2, 0
"00110000010000010000000001010100",	-- 8957: 	bgt	%r2, %r1, bgt_else.9250
"00111011110000010000000000000101",	-- 8958: 	lw	%r1, [%sp + 5]
"00111111111111100000000000000110",	-- 8959: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8960: 	addi	%sp, %sp, 7
"01011000000000000000011010101000",	-- 8961: 	jal	p_calc_diffuse.2670
"10101011110111100000000000000111",	-- 8962: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8963: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000100",	-- 8964: 	lw	%r2, [%sp + 4]
"10000100001000100000100000000000",	-- 8965: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 8966: 	lw	%r1, [%r1 + 0]
"11001100000000110000000000000000",	-- 8967: 	lli	%r3, 0
"00101000001000110000000000000010",	-- 8968: 	bneq	%r1, %r3, bneq_else.9251
"01010100000000000010001101001010",	-- 8969: 	j	bneq_cont.9252
	-- bneq_else.9251:
"00111011110000010000000000000101",	-- 8970: 	lw	%r1, [%sp + 5]
"00111111111111100000000000000110",	-- 8971: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8972: 	addi	%sp, %sp, 7
"01011000000000000000011010101110",	-- 8973: 	jal	p_group_id.2676
"10101011110111100000000000000111",	-- 8974: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8975: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000011",	-- 8976: 	lw	%r2, [%sp + 3]
"00111100001111100000000000000110",	-- 8977: 	sw	%r1, [%sp + 6]
"10000100000000100000100000000000",	-- 8978: 	add	%r1, %r0, %r2
"00111111111111100000000000000111",	-- 8979: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 8980: 	addi	%sp, %sp, 8
"01011000000000000000010100111000",	-- 8981: 	jal	vecbzero.2584
"10101011110111100000000000001000",	-- 8982: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8983: 	lw	%ra, [%sp + 7]
"00111011110000010000000000000101",	-- 8984: 	lw	%r1, [%sp + 5]
"00111111111111100000000000000111",	-- 8985: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 8986: 	addi	%sp, %sp, 8
"01011000000000000000011010111000",	-- 8987: 	jal	p_nvectors.2681
"10101011110111100000000000001000",	-- 8988: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8989: 	lw	%ra, [%sp + 7]
"00111011110000100000000000000101",	-- 8990: 	lw	%r2, [%sp + 5]
"00111100001111100000000000000111",	-- 8991: 	sw	%r1, [%sp + 7]
"10000100000000100000100000000000",	-- 8992: 	add	%r1, %r0, %r2
"00111111111111100000000000001000",	-- 8993: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 8994: 	addi	%sp, %sp, 9
"01011000000000000000011010100100",	-- 8995: 	jal	p_intersection_points.2666
"10101011110111100000000000001001",	-- 8996: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 8997: 	lw	%ra, [%sp + 8]
"00111011110000100000000000000110",	-- 8998: 	lw	%r2, [%sp + 6]
"00111011110000110000000000000010",	-- 8999: 	lw	%r3, [%sp + 2]
"10000100011000100001000000000000",	-- 9000: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 9001: 	lw	%r2, [%r2 + 0]
"00111011110000110000000000000100",	-- 9002: 	lw	%r3, [%sp + 4]
"00111011110001000000000000000111",	-- 9003: 	lw	%r4, [%sp + 7]
"10000100100000110010000000000000",	-- 9004: 	add	%r4, %r4, %r3
"00111000100001000000000000000000",	-- 9005: 	lw	%r4, [%r4 + 0]
"10000100001000110000100000000000",	-- 9006: 	add	%r1, %r1, %r3
"00111000001000010000000000000000",	-- 9007: 	lw	%r1, [%r1 + 0]
"00111011110110110000000000000001",	-- 9008: 	lw	%r27, [%sp + 1]
"10000100000000010001100000000000",	-- 9009: 	add	%r3, %r0, %r1
"10000100000000100000100000000000",	-- 9010: 	add	%r1, %r0, %r2
"10000100000001000001000000000000",	-- 9011: 	add	%r2, %r0, %r4
"00111111111111100000000000001000",	-- 9012: 	sw	%ra, [%sp + 8]
"00111011011110100000000000000000",	-- 9013: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001001",	-- 9014: 	addi	%sp, %sp, 9
"01010011010000000000000000000000",	-- 9015: 	jalr	%r26
"10101011110111100000000000001001",	-- 9016: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 9017: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000101",	-- 9018: 	lw	%r1, [%sp + 5]
"00111111111111100000000000001000",	-- 9019: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 9020: 	addi	%sp, %sp, 9
"01011000000000000000011010101100",	-- 9021: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000001001",	-- 9022: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 9023: 	lw	%ra, [%sp + 8]
"00111011110000100000000000000100",	-- 9024: 	lw	%r2, [%sp + 4]
"10000100001000100000100000000000",	-- 9025: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 9026: 	lw	%r1, [%r1 + 0]
"00111011110000110000000000000011",	-- 9027: 	lw	%r3, [%sp + 3]
"10000100000000110001000000000000",	-- 9028: 	add	%r2, %r0, %r3
"00111111111111100000000000001000",	-- 9029: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 9030: 	addi	%sp, %sp, 9
"01011000000000000000010100111011",	-- 9031: 	jal	veccpy.2586
"10101011110111100000000000001001",	-- 9032: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 9033: 	lw	%ra, [%sp + 8]
	-- bneq_cont.9252:
"11001100000000010000000000000001",	-- 9034: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 9035: 	lw	%r2, [%sp + 4]
"10000100010000010001000000000000",	-- 9036: 	add	%r2, %r2, %r1
"00111011110000010000000000000101",	-- 9037: 	lw	%r1, [%sp + 5]
"00111011110110110000000000000000",	-- 9038: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 9039: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 9040: 	jr	%r26
	-- bgt_else.9250:
"01001111111000000000000000000000",	-- 9041: 	jr	%ra
	-- bgt_else.9249:
"01001111111000000000000000000000",	-- 9042: 	jr	%ra
	-- pretrace_pixels.2966:
"00111011011001000000000000001001",	-- 9043: 	lw	%r4, [%r27 + 9]
"00111011011001010000000000001000",	-- 9044: 	lw	%r5, [%r27 + 8]
"00111011011001100000000000000111",	-- 9045: 	lw	%r6, [%r27 + 7]
"00111011011001110000000000000110",	-- 9046: 	lw	%r7, [%r27 + 6]
"00111011011010000000000000000101",	-- 9047: 	lw	%r8, [%r27 + 5]
"00111011011010010000000000000100",	-- 9048: 	lw	%r9, [%r27 + 4]
"00111011011010100000000000000011",	-- 9049: 	lw	%r10, [%r27 + 3]
"00111011011010110000000000000010",	-- 9050: 	lw	%r11, [%r27 + 2]
"00111011011011000000000000000001",	-- 9051: 	lw	%r12, [%r27 + 1]
"11001100000011010000000000000000",	-- 9052: 	lli	%r13, 0
"00110001101000100000000010100100",	-- 9053: 	bgt	%r13, %r2, bgt_else.9255
"11001100000011010000000000000000",	-- 9054: 	lli	%r13, 0
"10000101000011010100000000000000",	-- 9055: 	add	%r8, %r8, %r13
"10010001000000110000000000000000",	-- 9056: 	lf	%f3, [%r8 + 0]
"11001100000010000000000000000000",	-- 9057: 	lli	%r8, 0
"10000101100010000100000000000000",	-- 9058: 	add	%r8, %r12, %r8
"00111001000010000000000000000000",	-- 9059: 	lw	%r8, [%r8 + 0]
"10001000010010000100000000000000",	-- 9060: 	sub	%r8, %r2, %r8
"00111111011111100000000000000000",	-- 9061: 	sw	%r27, [%sp + 0]
"00111101011111100000000000000001",	-- 9062: 	sw	%r11, [%sp + 1]
"00111100011111100000000000000010",	-- 9063: 	sw	%r3, [%sp + 2]
"00111100101111100000000000000011",	-- 9064: 	sw	%r5, [%sp + 3]
"00111100010111100000000000000100",	-- 9065: 	sw	%r2, [%sp + 4]
"00111100001111100000000000000101",	-- 9066: 	sw	%r1, [%sp + 5]
"00111100100111100000000000000110",	-- 9067: 	sw	%r4, [%sp + 6]
"00111100110111100000000000000111",	-- 9068: 	sw	%r6, [%sp + 7]
"00111101001111100000000000001000",	-- 9069: 	sw	%r9, [%sp + 8]
"10110000010111100000000000001001",	-- 9070: 	sf	%f2, [%sp + 9]
"10110000001111100000000000001010",	-- 9071: 	sf	%f1, [%sp + 10]
"00111101010111100000000000001011",	-- 9072: 	sw	%r10, [%sp + 11]
"10110000000111100000000000001100",	-- 9073: 	sf	%f0, [%sp + 12]
"00111100111111100000000000001101",	-- 9074: 	sw	%r7, [%sp + 13]
"10110000011111100000000000001110",	-- 9075: 	sf	%f3, [%sp + 14]
"10000100000010000000100000000000",	-- 9076: 	add	%r1, %r0, %r8
"00111111111111100000000000001111",	-- 9077: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9078: 	addi	%sp, %sp, 16
"01011000000000000010101000101010",	-- 9079: 	jal	yj_float_of_int
"10101011110111100000000000010000",	-- 9080: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9081: 	lw	%ra, [%sp + 15]
"10010011110000010000000000001110",	-- 9082: 	lf	%f1, [%sp + 14]
"11101000001000000000000000000000",	-- 9083: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 9084: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 9085: 	lli	%r2, 0
"00111011110000110000000000001101",	-- 9086: 	lw	%r3, [%sp + 13]
"10000100011000100001000000000000",	-- 9087: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 9088: 	lf	%f1, [%r2 + 0]
"11101000000000010000100000000000",	-- 9089: 	mulf	%f1, %f0, %f1
"10010011110000100000000000001100",	-- 9090: 	lf	%f2, [%sp + 12]
"11100000001000100000100000000000",	-- 9091: 	addf	%f1, %f1, %f2
"00111011110000100000000000001011",	-- 9092: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 9093: 	add	%r1, %r2, %r1
"10110000001000010000000000000000",	-- 9094: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000001",	-- 9095: 	lli	%r1, 1
"11001100000001000000000000000001",	-- 9096: 	lli	%r4, 1
"10000100011001000010000000000000",	-- 9097: 	add	%r4, %r3, %r4
"10010000100000010000000000000000",	-- 9098: 	lf	%f1, [%r4 + 0]
"11101000000000010000100000000000",	-- 9099: 	mulf	%f1, %f0, %f1
"10010011110000110000000000001010",	-- 9100: 	lf	%f3, [%sp + 10]
"11100000001000110000100000000000",	-- 9101: 	addf	%f1, %f1, %f3
"10000100010000010000100000000000",	-- 9102: 	add	%r1, %r2, %r1
"10110000001000010000000000000000",	-- 9103: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 9104: 	lli	%r1, 2
"11001100000001000000000000000010",	-- 9105: 	lli	%r4, 2
"10000100011001000001100000000000",	-- 9106: 	add	%r3, %r3, %r4
"10010000011000010000000000000000",	-- 9107: 	lf	%f1, [%r3 + 0]
"11101000000000010000000000000000",	-- 9108: 	mulf	%f0, %f0, %f1
"10010011110000010000000000001001",	-- 9109: 	lf	%f1, [%sp + 9]
"11100000000000010000000000000000",	-- 9110: 	addf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 9111: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 9112: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 9113: 	lli	%r1, 0
"10000100000000101101000000000000",	-- 9114: 	add	%r26, %r0, %r2
"10000100000000010001000000000000",	-- 9115: 	add	%r2, %r0, %r1
"10000100000110100000100000000000",	-- 9116: 	add	%r1, %r0, %r26
"00111111111111100000000000001111",	-- 9117: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9118: 	addi	%sp, %sp, 16
"01011000000000000000010101001110",	-- 9119: 	jal	vecunit_sgn.2594
"10101011110111100000000000010000",	-- 9120: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9121: 	lw	%ra, [%sp + 15]
"00111011110000010000000000001000",	-- 9122: 	lw	%r1, [%sp + 8]
"00111111111111100000000000001111",	-- 9123: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9124: 	addi	%sp, %sp, 16
"01011000000000000000010100111000",	-- 9125: 	jal	vecbzero.2584
"10101011110111100000000000010000",	-- 9126: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9127: 	lw	%ra, [%sp + 15]
"00111011110000010000000000000111",	-- 9128: 	lw	%r1, [%sp + 7]
"00111011110000100000000000000110",	-- 9129: 	lw	%r2, [%sp + 6]
"00111111111111100000000000001111",	-- 9130: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9131: 	addi	%sp, %sp, 16
"01011000000000000000010100111011",	-- 9132: 	jal	veccpy.2586
"10101011110111100000000000010000",	-- 9133: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9134: 	lw	%ra, [%sp + 15]
"11001100000000010000000000000000",	-- 9135: 	lli	%r1, 0
"00010100000000000000000000000000",	-- 9136: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 9137: 	lhif	%f0, 1.000000
"00111011110000100000000000000100",	-- 9138: 	lw	%r2, [%sp + 4]
"00111011110000110000000000000101",	-- 9139: 	lw	%r3, [%sp + 5]
"10000100011000100010000000000000",	-- 9140: 	add	%r4, %r3, %r2
"00111000100001000000000000000000",	-- 9141: 	lw	%r4, [%r4 + 0]
"00010100000000010000000000000000",	-- 9142: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 9143: 	lhif	%f1, 0.000000
"00111011110001010000000000001011",	-- 9144: 	lw	%r5, [%sp + 11]
"00111011110110110000000000000011",	-- 9145: 	lw	%r27, [%sp + 3]
"10000100000001000001100000000000",	-- 9146: 	add	%r3, %r0, %r4
"10000100000001010001000000000000",	-- 9147: 	add	%r2, %r0, %r5
"00111111111111100000000000001111",	-- 9148: 	sw	%ra, [%sp + 15]
"00111011011110100000000000000000",	-- 9149: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010000",	-- 9150: 	addi	%sp, %sp, 16
"01010011010000000000000000000000",	-- 9151: 	jalr	%r26
"10101011110111100000000000010000",	-- 9152: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9153: 	lw	%ra, [%sp + 15]
"00111011110000010000000000000100",	-- 9154: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000101",	-- 9155: 	lw	%r2, [%sp + 5]
"10000100010000010001100000000000",	-- 9156: 	add	%r3, %r2, %r1
"00111000011000110000000000000000",	-- 9157: 	lw	%r3, [%r3 + 0]
"10000100000000110000100000000000",	-- 9158: 	add	%r1, %r0, %r3
"00111111111111100000000000001111",	-- 9159: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9160: 	addi	%sp, %sp, 16
"01011000000000000000011010100010",	-- 9161: 	jal	p_rgb.2664
"10101011110111100000000000010000",	-- 9162: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9163: 	lw	%ra, [%sp + 15]
"00111011110000100000000000001000",	-- 9164: 	lw	%r2, [%sp + 8]
"00111111111111100000000000001111",	-- 9165: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9166: 	addi	%sp, %sp, 16
"01011000000000000000010100111011",	-- 9167: 	jal	veccpy.2586
"10101011110111100000000000010000",	-- 9168: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9169: 	lw	%ra, [%sp + 15]
"00111011110000010000000000000100",	-- 9170: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000101",	-- 9171: 	lw	%r2, [%sp + 5]
"10000100010000010001100000000000",	-- 9172: 	add	%r3, %r2, %r1
"00111000011000110000000000000000",	-- 9173: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000000010",	-- 9174: 	lw	%r4, [%sp + 2]
"10000100000001000001000000000000",	-- 9175: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 9176: 	add	%r1, %r0, %r3
"00111111111111100000000000001111",	-- 9177: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9178: 	addi	%sp, %sp, 16
"01011000000000000000011010110011",	-- 9179: 	jal	p_set_group_id.2678
"10101011110111100000000000010000",	-- 9180: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9181: 	lw	%ra, [%sp + 15]
"00111011110000010000000000000100",	-- 9182: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000101",	-- 9183: 	lw	%r2, [%sp + 5]
"10000100010000010001100000000000",	-- 9184: 	add	%r3, %r2, %r1
"00111000011000110000000000000000",	-- 9185: 	lw	%r3, [%r3 + 0]
"11001100000001000000000000000000",	-- 9186: 	lli	%r4, 0
"00111011110110110000000000000001",	-- 9187: 	lw	%r27, [%sp + 1]
"10000100000001000001000000000000",	-- 9188: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 9189: 	add	%r1, %r0, %r3
"00111111111111100000000000001111",	-- 9190: 	sw	%ra, [%sp + 15]
"00111011011110100000000000000000",	-- 9191: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010000",	-- 9192: 	addi	%sp, %sp, 16
"01010011010000000000000000000000",	-- 9193: 	jalr	%r26
"10101011110111100000000000010000",	-- 9194: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9195: 	lw	%ra, [%sp + 15]
"11001100000000010000000000000001",	-- 9196: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 9197: 	lw	%r2, [%sp + 4]
"10001000010000010000100000000000",	-- 9198: 	sub	%r1, %r2, %r1
"11001100000000100000000000000001",	-- 9199: 	lli	%r2, 1
"00111011110000110000000000000010",	-- 9200: 	lw	%r3, [%sp + 2]
"00111100001111100000000000001111",	-- 9201: 	sw	%r1, [%sp + 15]
"10000100000000110000100000000000",	-- 9202: 	add	%r1, %r0, %r3
"00111111111111100000000000010000",	-- 9203: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 9204: 	addi	%sp, %sp, 17
"01011000000000000000010100011101",	-- 9205: 	jal	add_mod5.2573
"10101011110111100000000000010001",	-- 9206: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 9207: 	lw	%ra, [%sp + 16]
"10000100000000010001100000000000",	-- 9208: 	add	%r3, %r0, %r1
"10010011110000000000000000001100",	-- 9209: 	lf	%f0, [%sp + 12]
"10010011110000010000000000001010",	-- 9210: 	lf	%f1, [%sp + 10]
"10010011110000100000000000001001",	-- 9211: 	lf	%f2, [%sp + 9]
"00111011110000010000000000000101",	-- 9212: 	lw	%r1, [%sp + 5]
"00111011110000100000000000001111",	-- 9213: 	lw	%r2, [%sp + 15]
"00111011110110110000000000000000",	-- 9214: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 9215: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 9216: 	jr	%r26
	-- bgt_else.9255:
"01001111111000000000000000000000",	-- 9217: 	jr	%ra
	-- pretrace_line.2973:
"00111011011001000000000000000110",	-- 9218: 	lw	%r4, [%r27 + 6]
"00111011011001010000000000000101",	-- 9219: 	lw	%r5, [%r27 + 5]
"00111011011001100000000000000100",	-- 9220: 	lw	%r6, [%r27 + 4]
"00111011011001110000000000000011",	-- 9221: 	lw	%r7, [%r27 + 3]
"00111011011010000000000000000010",	-- 9222: 	lw	%r8, [%r27 + 2]
"00111011011010010000000000000001",	-- 9223: 	lw	%r9, [%r27 + 1]
"11001100000010100000000000000000",	-- 9224: 	lli	%r10, 0
"10000100110010100011000000000000",	-- 9225: 	add	%r6, %r6, %r10
"10010000110000000000000000000000",	-- 9226: 	lf	%f0, [%r6 + 0]
"11001100000001100000000000000001",	-- 9227: 	lli	%r6, 1
"10000101001001100011000000000000",	-- 9228: 	add	%r6, %r9, %r6
"00111000110001100000000000000000",	-- 9229: 	lw	%r6, [%r6 + 0]
"10001000010001100001000000000000",	-- 9230: 	sub	%r2, %r2, %r6
"00111100011111100000000000000000",	-- 9231: 	sw	%r3, [%sp + 0]
"00111100001111100000000000000001",	-- 9232: 	sw	%r1, [%sp + 1]
"00111100111111100000000000000010",	-- 9233: 	sw	%r7, [%sp + 2]
"00111101000111100000000000000011",	-- 9234: 	sw	%r8, [%sp + 3]
"00111100100111100000000000000100",	-- 9235: 	sw	%r4, [%sp + 4]
"00111100101111100000000000000101",	-- 9236: 	sw	%r5, [%sp + 5]
"10110000000111100000000000000110",	-- 9237: 	sf	%f0, [%sp + 6]
"10000100000000100000100000000000",	-- 9238: 	add	%r1, %r0, %r2
"00111111111111100000000000000111",	-- 9239: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 9240: 	addi	%sp, %sp, 8
"01011000000000000010101000101010",	-- 9241: 	jal	yj_float_of_int
"10101011110111100000000000001000",	-- 9242: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 9243: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000110",	-- 9244: 	lf	%f1, [%sp + 6]
"11101000001000000000000000000000",	-- 9245: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 9246: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 9247: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 9248: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 9249: 	lf	%f1, [%r1 + 0]
"11101000000000010000100000000000",	-- 9250: 	mulf	%f1, %f0, %f1
"11001100000000010000000000000000",	-- 9251: 	lli	%r1, 0
"00111011110000110000000000000100",	-- 9252: 	lw	%r3, [%sp + 4]
"10000100011000010000100000000000",	-- 9253: 	add	%r1, %r3, %r1
"10010000001000100000000000000000",	-- 9254: 	lf	%f2, [%r1 + 0]
"11100000001000100000100000000000",	-- 9255: 	addf	%f1, %f1, %f2
"11001100000000010000000000000001",	-- 9256: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 9257: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 9258: 	lf	%f2, [%r1 + 0]
"11101000000000100001000000000000",	-- 9259: 	mulf	%f2, %f0, %f2
"11001100000000010000000000000001",	-- 9260: 	lli	%r1, 1
"10000100011000010000100000000000",	-- 9261: 	add	%r1, %r3, %r1
"10010000001000110000000000000000",	-- 9262: 	lf	%f3, [%r1 + 0]
"11100000010000110001000000000000",	-- 9263: 	addf	%f2, %f2, %f3
"11001100000000010000000000000010",	-- 9264: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 9265: 	add	%r1, %r2, %r1
"10010000001000110000000000000000",	-- 9266: 	lf	%f3, [%r1 + 0]
"11101000000000110000000000000000",	-- 9267: 	mulf	%f0, %f0, %f3
"11001100000000010000000000000010",	-- 9268: 	lli	%r1, 2
"10000100011000010000100000000000",	-- 9269: 	add	%r1, %r3, %r1
"10010000001000110000000000000000",	-- 9270: 	lf	%f3, [%r1 + 0]
"11100000000000110000000000000000",	-- 9271: 	addf	%f0, %f0, %f3
"11001100000000010000000000000000",	-- 9272: 	lli	%r1, 0
"00111011110000100000000000000011",	-- 9273: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 9274: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 9275: 	lw	%r1, [%r1 + 0]
"11001100000000100000000000000001",	-- 9276: 	lli	%r2, 1
"10001000001000100001000000000000",	-- 9277: 	sub	%r2, %r1, %r2
"00111011110000010000000000000001",	-- 9278: 	lw	%r1, [%sp + 1]
"00111011110000110000000000000000",	-- 9279: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000010",	-- 9280: 	lw	%r27, [%sp + 2]
"00001100010111110000000000000000",	-- 9281: 	movf	%f31, %f2
"00001100000000100000000000000000",	-- 9282: 	movf	%f2, %f0
"00001100001000000000000000000000",	-- 9283: 	movf	%f0, %f1
"00001111111000010000000000000000",	-- 9284: 	movf	%f1, %f31
"00111011011110100000000000000000",	-- 9285: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 9286: 	jr	%r26
	-- scan_pixel.2977:
"00111011011001100000000000000110",	-- 9287: 	lw	%r6, [%r27 + 6]
"00111011011001110000000000000101",	-- 9288: 	lw	%r7, [%r27 + 5]
"00111011011010000000000000000100",	-- 9289: 	lw	%r8, [%r27 + 4]
"00111011011010010000000000000011",	-- 9290: 	lw	%r9, [%r27 + 3]
"00111011011010100000000000000010",	-- 9291: 	lw	%r10, [%r27 + 2]
"00111011011010110000000000000001",	-- 9292: 	lw	%r11, [%r27 + 1]
"11001100000011000000000000000000",	-- 9293: 	lli	%r12, 0
"10000101010011000101000000000000",	-- 9294: 	add	%r10, %r10, %r12
"00111001010010100000000000000000",	-- 9295: 	lw	%r10, [%r10 + 0]
"00110001010000010000000000000010",	-- 9296: 	bgt	%r10, %r1, bgt_else.9257
"01001111111000000000000000000000",	-- 9297: 	jr	%ra
	-- bgt_else.9257:
"10000100100000010101000000000000",	-- 9298: 	add	%r10, %r4, %r1
"00111001010010100000000000000000",	-- 9299: 	lw	%r10, [%r10 + 0]
"00111111011111100000000000000000",	-- 9300: 	sw	%r27, [%sp + 0]
"00111100110111100000000000000001",	-- 9301: 	sw	%r6, [%sp + 1]
"00111100011111100000000000000010",	-- 9302: 	sw	%r3, [%sp + 2]
"00111100111111100000000000000011",	-- 9303: 	sw	%r7, [%sp + 3]
"00111101011111100000000000000100",	-- 9304: 	sw	%r11, [%sp + 4]
"00111100100111100000000000000101",	-- 9305: 	sw	%r4, [%sp + 5]
"00111100101111100000000000000110",	-- 9306: 	sw	%r5, [%sp + 6]
"00111100010111100000000000000111",	-- 9307: 	sw	%r2, [%sp + 7]
"00111100001111100000000000001000",	-- 9308: 	sw	%r1, [%sp + 8]
"00111101001111100000000000001001",	-- 9309: 	sw	%r9, [%sp + 9]
"00111101000111100000000000001010",	-- 9310: 	sw	%r8, [%sp + 10]
"10000100000010100000100000000000",	-- 9311: 	add	%r1, %r0, %r10
"00111111111111100000000000001011",	-- 9312: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 9313: 	addi	%sp, %sp, 12
"01011000000000000000011010100010",	-- 9314: 	jal	p_rgb.2664
"10101011110111100000000000001100",	-- 9315: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9316: 	lw	%ra, [%sp + 11]
"10000100000000010001000000000000",	-- 9317: 	add	%r2, %r0, %r1
"00111011110000010000000000001010",	-- 9318: 	lw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 9319: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 9320: 	addi	%sp, %sp, 12
"01011000000000000000010100111011",	-- 9321: 	jal	veccpy.2586
"10101011110111100000000000001100",	-- 9322: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9323: 	lw	%ra, [%sp + 11]
"00111011110000010000000000001000",	-- 9324: 	lw	%r1, [%sp + 8]
"00111011110000100000000000000111",	-- 9325: 	lw	%r2, [%sp + 7]
"00111011110000110000000000000110",	-- 9326: 	lw	%r3, [%sp + 6]
"00111011110110110000000000001001",	-- 9327: 	lw	%r27, [%sp + 9]
"00111111111111100000000000001011",	-- 9328: 	sw	%ra, [%sp + 11]
"00111011011110100000000000000000",	-- 9329: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001100",	-- 9330: 	addi	%sp, %sp, 12
"01010011010000000000000000000000",	-- 9331: 	jalr	%r26
"10101011110111100000000000001100",	-- 9332: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9333: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 9334: 	lli	%r2, 0
"00101000001000100000000000010000",	-- 9335: 	bneq	%r1, %r2, bneq_else.9259
"00111011110000010000000000001000",	-- 9336: 	lw	%r1, [%sp + 8]
"00111011110000100000000000000101",	-- 9337: 	lw	%r2, [%sp + 5]
"10000100010000010001100000000000",	-- 9338: 	add	%r3, %r2, %r1
"00111000011000110000000000000000",	-- 9339: 	lw	%r3, [%r3 + 0]
"11001100000001000000000000000000",	-- 9340: 	lli	%r4, 0
"00111011110110110000000000000100",	-- 9341: 	lw	%r27, [%sp + 4]
"10000100000001000001000000000000",	-- 9342: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 9343: 	add	%r1, %r0, %r3
"00111111111111100000000000001011",	-- 9344: 	sw	%ra, [%sp + 11]
"00111011011110100000000000000000",	-- 9345: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001100",	-- 9346: 	addi	%sp, %sp, 12
"01010011010000000000000000000000",	-- 9347: 	jalr	%r26
"10101011110111100000000000001100",	-- 9348: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9349: 	lw	%ra, [%sp + 11]
"01010100000000000010010010010100",	-- 9350: 	j	bneq_cont.9260
	-- bneq_else.9259:
"11001100000001100000000000000000",	-- 9351: 	lli	%r6, 0
"00111011110000010000000000001000",	-- 9352: 	lw	%r1, [%sp + 8]
"00111011110000100000000000000111",	-- 9353: 	lw	%r2, [%sp + 7]
"00111011110000110000000000000010",	-- 9354: 	lw	%r3, [%sp + 2]
"00111011110001000000000000000101",	-- 9355: 	lw	%r4, [%sp + 5]
"00111011110001010000000000000110",	-- 9356: 	lw	%r5, [%sp + 6]
"00111011110110110000000000000011",	-- 9357: 	lw	%r27, [%sp + 3]
"00111111111111100000000000001011",	-- 9358: 	sw	%ra, [%sp + 11]
"00111011011110100000000000000000",	-- 9359: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001100",	-- 9360: 	addi	%sp, %sp, 12
"01010011010000000000000000000000",	-- 9361: 	jalr	%r26
"10101011110111100000000000001100",	-- 9362: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9363: 	lw	%ra, [%sp + 11]
	-- bneq_cont.9260:
"00111011110110110000000000000001",	-- 9364: 	lw	%r27, [%sp + 1]
"00111111111111100000000000001011",	-- 9365: 	sw	%ra, [%sp + 11]
"00111011011110100000000000000000",	-- 9366: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001100",	-- 9367: 	addi	%sp, %sp, 12
"01010011010000000000000000000000",	-- 9368: 	jalr	%r26
"10101011110111100000000000001100",	-- 9369: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9370: 	lw	%ra, [%sp + 11]
"11001100000000010000000000000001",	-- 9371: 	lli	%r1, 1
"00111011110000100000000000001000",	-- 9372: 	lw	%r2, [%sp + 8]
"10000100010000010000100000000000",	-- 9373: 	add	%r1, %r2, %r1
"00111011110000100000000000000111",	-- 9374: 	lw	%r2, [%sp + 7]
"00111011110000110000000000000010",	-- 9375: 	lw	%r3, [%sp + 2]
"00111011110001000000000000000101",	-- 9376: 	lw	%r4, [%sp + 5]
"00111011110001010000000000000110",	-- 9377: 	lw	%r5, [%sp + 6]
"00111011110110110000000000000000",	-- 9378: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 9379: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 9380: 	jr	%r26
	-- scan_line.2983:
"00111011011001100000000000000011",	-- 9381: 	lw	%r6, [%r27 + 3]
"00111011011001110000000000000010",	-- 9382: 	lw	%r7, [%r27 + 2]
"00111011011010000000000000000001",	-- 9383: 	lw	%r8, [%r27 + 1]
"11001100000010010000000000000001",	-- 9384: 	lli	%r9, 1
"10000101000010010100100000000000",	-- 9385: 	add	%r9, %r8, %r9
"00111001001010010000000000000000",	-- 9386: 	lw	%r9, [%r9 + 0]
"00110001001000010000000000000010",	-- 9387: 	bgt	%r9, %r1, bgt_else.9261
"01001111111000000000000000000000",	-- 9388: 	jr	%ra
	-- bgt_else.9261:
"11001100000010010000000000000001",	-- 9389: 	lli	%r9, 1
"10000101000010010100000000000000",	-- 9390: 	add	%r8, %r8, %r9
"00111001000010000000000000000000",	-- 9391: 	lw	%r8, [%r8 + 0]
"11001100000010010000000000000001",	-- 9392: 	lli	%r9, 1
"10001001000010010100000000000000",	-- 9393: 	sub	%r8, %r8, %r9
"00111111011111100000000000000000",	-- 9394: 	sw	%r27, [%sp + 0]
"00111100101111100000000000000001",	-- 9395: 	sw	%r5, [%sp + 1]
"00111100100111100000000000000010",	-- 9396: 	sw	%r4, [%sp + 2]
"00111100011111100000000000000011",	-- 9397: 	sw	%r3, [%sp + 3]
"00111100010111100000000000000100",	-- 9398: 	sw	%r2, [%sp + 4]
"00111100001111100000000000000101",	-- 9399: 	sw	%r1, [%sp + 5]
"00111100110111100000000000000110",	-- 9400: 	sw	%r6, [%sp + 6]
"00110001000000010000000000000010",	-- 9401: 	bgt	%r8, %r1, bgt_else.9263
"01010100000000000010010011000111",	-- 9402: 	j	bgt_cont.9264
	-- bgt_else.9263:
"11001100000010000000000000000001",	-- 9403: 	lli	%r8, 1
"10000100001010000100000000000000",	-- 9404: 	add	%r8, %r1, %r8
"10000100000001010001100000000000",	-- 9405: 	add	%r3, %r0, %r5
"10000100000010000001000000000000",	-- 9406: 	add	%r2, %r0, %r8
"10000100000001000000100000000000",	-- 9407: 	add	%r1, %r0, %r4
"10000100000001111101100000000000",	-- 9408: 	add	%r27, %r0, %r7
"00111111111111100000000000000111",	-- 9409: 	sw	%ra, [%sp + 7]
"00111011011110100000000000000000",	-- 9410: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001000",	-- 9411: 	addi	%sp, %sp, 8
"01010011010000000000000000000000",	-- 9412: 	jalr	%r26
"10101011110111100000000000001000",	-- 9413: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 9414: 	lw	%ra, [%sp + 7]
	-- bgt_cont.9264:
"11001100000000010000000000000000",	-- 9415: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 9416: 	lw	%r2, [%sp + 5]
"00111011110000110000000000000100",	-- 9417: 	lw	%r3, [%sp + 4]
"00111011110001000000000000000011",	-- 9418: 	lw	%r4, [%sp + 3]
"00111011110001010000000000000010",	-- 9419: 	lw	%r5, [%sp + 2]
"00111011110110110000000000000110",	-- 9420: 	lw	%r27, [%sp + 6]
"00111111111111100000000000000111",	-- 9421: 	sw	%ra, [%sp + 7]
"00111011011110100000000000000000",	-- 9422: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001000",	-- 9423: 	addi	%sp, %sp, 8
"01010011010000000000000000000000",	-- 9424: 	jalr	%r26
"10101011110111100000000000001000",	-- 9425: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 9426: 	lw	%ra, [%sp + 7]
"11001100000000010000000000000001",	-- 9427: 	lli	%r1, 1
"00111011110000100000000000000101",	-- 9428: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 9429: 	add	%r1, %r2, %r1
"11001100000000100000000000000010",	-- 9430: 	lli	%r2, 2
"00111011110000110000000000000001",	-- 9431: 	lw	%r3, [%sp + 1]
"00111100001111100000000000000111",	-- 9432: 	sw	%r1, [%sp + 7]
"10000100000000110000100000000000",	-- 9433: 	add	%r1, %r0, %r3
"00111111111111100000000000001000",	-- 9434: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 9435: 	addi	%sp, %sp, 9
"01011000000000000000010100011101",	-- 9436: 	jal	add_mod5.2573
"10101011110111100000000000001001",	-- 9437: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 9438: 	lw	%ra, [%sp + 8]
"10000100000000010010100000000000",	-- 9439: 	add	%r5, %r0, %r1
"00111011110000010000000000000111",	-- 9440: 	lw	%r1, [%sp + 7]
"00111011110000100000000000000011",	-- 9441: 	lw	%r2, [%sp + 3]
"00111011110000110000000000000010",	-- 9442: 	lw	%r3, [%sp + 2]
"00111011110001000000000000000100",	-- 9443: 	lw	%r4, [%sp + 4]
"00111011110110110000000000000000",	-- 9444: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 9445: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 9446: 	jr	%r26
	-- create_float5x3array.2989:
"11001100000000010000000000000011",	-- 9447: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 9448: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9449: 	lhif	%f0, 0.000000
"00111111111111100000000000000000",	-- 9450: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 9451: 	addi	%sp, %sp, 1
"01011000000000000010101000100010",	-- 9452: 	jal	yj_create_float_array
"10101011110111100000000000000001",	-- 9453: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 9454: 	lw	%ra, [%sp + 0]
"10000100000000010001000000000000",	-- 9455: 	add	%r2, %r0, %r1
"11001100000000010000000000000101",	-- 9456: 	lli	%r1, 5
"00111111111111100000000000000000",	-- 9457: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 9458: 	addi	%sp, %sp, 1
"01011000000000000010101000011010",	-- 9459: 	jal	yj_create_array
"10101011110111100000000000000001",	-- 9460: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 9461: 	lw	%ra, [%sp + 0]
"11001100000000100000000000000001",	-- 9462: 	lli	%r2, 1
"11001100000000110000000000000011",	-- 9463: 	lli	%r3, 3
"00010100000000000000000000000000",	-- 9464: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9465: 	lhif	%f0, 0.000000
"00111100010111100000000000000000",	-- 9466: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 9467: 	sw	%r1, [%sp + 1]
"10000100000000110000100000000000",	-- 9468: 	add	%r1, %r0, %r3
"00111111111111100000000000000010",	-- 9469: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9470: 	addi	%sp, %sp, 3
"01011000000000000010101000100010",	-- 9471: 	jal	yj_create_float_array
"10101011110111100000000000000011",	-- 9472: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9473: 	lw	%ra, [%sp + 2]
"00111011110000100000000000000000",	-- 9474: 	lw	%r2, [%sp + 0]
"00111011110000110000000000000001",	-- 9475: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 9476: 	add	%r2, %r3, %r2
"00111100001000100000000000000000",	-- 9477: 	sw	%r1, [%r2 + 0]
"11001100000000010000000000000010",	-- 9478: 	lli	%r1, 2
"11001100000000100000000000000011",	-- 9479: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 9480: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9481: 	lhif	%f0, 0.000000
"00111100001111100000000000000010",	-- 9482: 	sw	%r1, [%sp + 2]
"10000100000000100000100000000000",	-- 9483: 	add	%r1, %r0, %r2
"00111111111111100000000000000011",	-- 9484: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 9485: 	addi	%sp, %sp, 4
"01011000000000000010101000100010",	-- 9486: 	jal	yj_create_float_array
"10101011110111100000000000000100",	-- 9487: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 9488: 	lw	%ra, [%sp + 3]
"00111011110000100000000000000010",	-- 9489: 	lw	%r2, [%sp + 2]
"00111011110000110000000000000001",	-- 9490: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 9491: 	add	%r2, %r3, %r2
"00111100001000100000000000000000",	-- 9492: 	sw	%r1, [%r2 + 0]
"11001100000000010000000000000011",	-- 9493: 	lli	%r1, 3
"11001100000000100000000000000011",	-- 9494: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 9495: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9496: 	lhif	%f0, 0.000000
"00111100001111100000000000000011",	-- 9497: 	sw	%r1, [%sp + 3]
"10000100000000100000100000000000",	-- 9498: 	add	%r1, %r0, %r2
"00111111111111100000000000000100",	-- 9499: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 9500: 	addi	%sp, %sp, 5
"01011000000000000010101000100010",	-- 9501: 	jal	yj_create_float_array
"10101011110111100000000000000101",	-- 9502: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 9503: 	lw	%ra, [%sp + 4]
"00111011110000100000000000000011",	-- 9504: 	lw	%r2, [%sp + 3]
"00111011110000110000000000000001",	-- 9505: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 9506: 	add	%r2, %r3, %r2
"00111100001000100000000000000000",	-- 9507: 	sw	%r1, [%r2 + 0]
"11001100000000010000000000000100",	-- 9508: 	lli	%r1, 4
"11001100000000100000000000000011",	-- 9509: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 9510: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9511: 	lhif	%f0, 0.000000
"00111100001111100000000000000100",	-- 9512: 	sw	%r1, [%sp + 4]
"10000100000000100000100000000000",	-- 9513: 	add	%r1, %r0, %r2
"00111111111111100000000000000101",	-- 9514: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 9515: 	addi	%sp, %sp, 6
"01011000000000000010101000100010",	-- 9516: 	jal	yj_create_float_array
"10101011110111100000000000000110",	-- 9517: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 9518: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000100",	-- 9519: 	lw	%r2, [%sp + 4]
"00111011110000110000000000000001",	-- 9520: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 9521: 	add	%r2, %r3, %r2
"00111100001000100000000000000000",	-- 9522: 	sw	%r1, [%r2 + 0]
"10000100000000110000100000000000",	-- 9523: 	add	%r1, %r0, %r3
"01001111111000000000000000000000",	-- 9524: 	jr	%ra
	-- create_pixel.2991:
"11001100000000010000000000000011",	-- 9525: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 9526: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9527: 	lhif	%f0, 0.000000
"00111111111111100000000000000000",	-- 9528: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 9529: 	addi	%sp, %sp, 1
"01011000000000000010101000100010",	-- 9530: 	jal	yj_create_float_array
"10101011110111100000000000000001",	-- 9531: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 9532: 	lw	%ra, [%sp + 0]
"00111100001111100000000000000000",	-- 9533: 	sw	%r1, [%sp + 0]
"00111111111111100000000000000001",	-- 9534: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 9535: 	addi	%sp, %sp, 2
"01011000000000000010010011100111",	-- 9536: 	jal	create_float5x3array.2989
"10101011110111100000000000000010",	-- 9537: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 9538: 	lw	%ra, [%sp + 1]
"11001100000000100000000000000101",	-- 9539: 	lli	%r2, 5
"11001100000000110000000000000000",	-- 9540: 	lli	%r3, 0
"00111100001111100000000000000001",	-- 9541: 	sw	%r1, [%sp + 1]
"10000100000000100000100000000000",	-- 9542: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 9543: 	add	%r2, %r0, %r3
"00111111111111100000000000000010",	-- 9544: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9545: 	addi	%sp, %sp, 3
"01011000000000000010101000011010",	-- 9546: 	jal	yj_create_array
"10101011110111100000000000000011",	-- 9547: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9548: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000101",	-- 9549: 	lli	%r2, 5
"11001100000000110000000000000000",	-- 9550: 	lli	%r3, 0
"00111100001111100000000000000010",	-- 9551: 	sw	%r1, [%sp + 2]
"10000100000000100000100000000000",	-- 9552: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 9553: 	add	%r2, %r0, %r3
"00111111111111100000000000000011",	-- 9554: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 9555: 	addi	%sp, %sp, 4
"01011000000000000010101000011010",	-- 9556: 	jal	yj_create_array
"10101011110111100000000000000100",	-- 9557: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 9558: 	lw	%ra, [%sp + 3]
"00111100001111100000000000000011",	-- 9559: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 9560: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 9561: 	addi	%sp, %sp, 5
"01011000000000000010010011100111",	-- 9562: 	jal	create_float5x3array.2989
"10101011110111100000000000000101",	-- 9563: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 9564: 	lw	%ra, [%sp + 4]
"00111100001111100000000000000100",	-- 9565: 	sw	%r1, [%sp + 4]
"00111111111111100000000000000101",	-- 9566: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 9567: 	addi	%sp, %sp, 6
"01011000000000000010010011100111",	-- 9568: 	jal	create_float5x3array.2989
"10101011110111100000000000000110",	-- 9569: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 9570: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000001",	-- 9571: 	lli	%r2, 1
"11001100000000110000000000000000",	-- 9572: 	lli	%r3, 0
"00111100001111100000000000000101",	-- 9573: 	sw	%r1, [%sp + 5]
"10000100000000100000100000000000",	-- 9574: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 9575: 	add	%r2, %r0, %r3
"00111111111111100000000000000110",	-- 9576: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 9577: 	addi	%sp, %sp, 7
"01011000000000000010101000011010",	-- 9578: 	jal	yj_create_array
"10101011110111100000000000000111",	-- 9579: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 9580: 	lw	%ra, [%sp + 6]
"00111100001111100000000000000110",	-- 9581: 	sw	%r1, [%sp + 6]
"00111111111111100000000000000111",	-- 9582: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 9583: 	addi	%sp, %sp, 8
"01011000000000000010010011100111",	-- 9584: 	jal	create_float5x3array.2989
"10101011110111100000000000001000",	-- 9585: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 9586: 	lw	%ra, [%sp + 7]
"10000100000111010001000000000000",	-- 9587: 	add	%r2, %r0, %hp
"10100111101111010000000000001000",	-- 9588: 	addi	%hp, %hp, 8
"00111100001000100000000000000111",	-- 9589: 	sw	%r1, [%r2 + 7]
"00111011110000010000000000000110",	-- 9590: 	lw	%r1, [%sp + 6]
"00111100001000100000000000000110",	-- 9591: 	sw	%r1, [%r2 + 6]
"00111011110000010000000000000101",	-- 9592: 	lw	%r1, [%sp + 5]
"00111100001000100000000000000101",	-- 9593: 	sw	%r1, [%r2 + 5]
"00111011110000010000000000000100",	-- 9594: 	lw	%r1, [%sp + 4]
"00111100001000100000000000000100",	-- 9595: 	sw	%r1, [%r2 + 4]
"00111011110000010000000000000011",	-- 9596: 	lw	%r1, [%sp + 3]
"00111100001000100000000000000011",	-- 9597: 	sw	%r1, [%r2 + 3]
"00111011110000010000000000000010",	-- 9598: 	lw	%r1, [%sp + 2]
"00111100001000100000000000000010",	-- 9599: 	sw	%r1, [%r2 + 2]
"00111011110000010000000000000001",	-- 9600: 	lw	%r1, [%sp + 1]
"00111100001000100000000000000001",	-- 9601: 	sw	%r1, [%r2 + 1]
"00111011110000010000000000000000",	-- 9602: 	lw	%r1, [%sp + 0]
"00111100001000100000000000000000",	-- 9603: 	sw	%r1, [%r2 + 0]
"10000100000000100000100000000000",	-- 9604: 	add	%r1, %r0, %r2
"01001111111000000000000000000000",	-- 9605: 	jr	%ra
	-- init_line_elements.2993:
"11001100000000110000000000000000",	-- 9606: 	lli	%r3, 0
"00110000011000100000000000010000",	-- 9607: 	bgt	%r3, %r2, bgt_else.9265
"00111100010111100000000000000000",	-- 9608: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 9609: 	sw	%r1, [%sp + 1]
"00111111111111100000000000000010",	-- 9610: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9611: 	addi	%sp, %sp, 3
"01011000000000000010010100110101",	-- 9612: 	jal	create_pixel.2991
"10101011110111100000000000000011",	-- 9613: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9614: 	lw	%ra, [%sp + 2]
"00111011110000100000000000000000",	-- 9615: 	lw	%r2, [%sp + 0]
"00111011110000110000000000000001",	-- 9616: 	lw	%r3, [%sp + 1]
"10000100011000100010000000000000",	-- 9617: 	add	%r4, %r3, %r2
"00111100001001000000000000000000",	-- 9618: 	sw	%r1, [%r4 + 0]
"11001100000000010000000000000001",	-- 9619: 	lli	%r1, 1
"10001000010000010001000000000000",	-- 9620: 	sub	%r2, %r2, %r1
"10000100000000110000100000000000",	-- 9621: 	add	%r1, %r0, %r3
"01010100000000000010010110000110",	-- 9622: 	j	init_line_elements.2993
	-- bgt_else.9265:
"01001111111000000000000000000000",	-- 9623: 	jr	%ra
	-- create_pixelline.2996:
"00111011011000010000000000000001",	-- 9624: 	lw	%r1, [%r27 + 1]
"11001100000000100000000000000000",	-- 9625: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 9626: 	add	%r2, %r1, %r2
"00111000010000100000000000000000",	-- 9627: 	lw	%r2, [%r2 + 0]
"00111100001111100000000000000000",	-- 9628: 	sw	%r1, [%sp + 0]
"00111100010111100000000000000001",	-- 9629: 	sw	%r2, [%sp + 1]
"00111111111111100000000000000010",	-- 9630: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9631: 	addi	%sp, %sp, 3
"01011000000000000010010100110101",	-- 9632: 	jal	create_pixel.2991
"10101011110111100000000000000011",	-- 9633: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9634: 	lw	%ra, [%sp + 2]
"10000100000000010001000000000000",	-- 9635: 	add	%r2, %r0, %r1
"00111011110000010000000000000001",	-- 9636: 	lw	%r1, [%sp + 1]
"00111111111111100000000000000010",	-- 9637: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9638: 	addi	%sp, %sp, 3
"01011000000000000010101000011010",	-- 9639: 	jal	yj_create_array
"10101011110111100000000000000011",	-- 9640: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9641: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000000",	-- 9642: 	lli	%r2, 0
"00111011110000110000000000000000",	-- 9643: 	lw	%r3, [%sp + 0]
"10000100011000100001000000000000",	-- 9644: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 9645: 	lw	%r2, [%r2 + 0]
"11001100000000110000000000000010",	-- 9646: 	lli	%r3, 2
"10001000010000110001000000000000",	-- 9647: 	sub	%r2, %r2, %r3
"01010100000000000010010110000110",	-- 9648: 	j	init_line_elements.2993
	-- tan.2998:
"10110000000111100000000000000000",	-- 9649: 	sf	%f0, [%sp + 0]
"00111111111111100000000000000001",	-- 9650: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 9651: 	addi	%sp, %sp, 2
"01011000000000000000010001010111",	-- 9652: 	jal	sin.2516
"10101011110111100000000000000010",	-- 9653: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 9654: 	lw	%ra, [%sp + 1]
"10010011110000010000000000000000",	-- 9655: 	lf	%f1, [%sp + 0]
"10110000000111100000000000000001",	-- 9656: 	sf	%f0, [%sp + 1]
"00001100001000000000000000000000",	-- 9657: 	movf	%f0, %f1
"00111111111111100000000000000010",	-- 9658: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9659: 	addi	%sp, %sp, 3
"01011000000000000000010010010110",	-- 9660: 	jal	cos.2518
"10101011110111100000000000000011",	-- 9661: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9662: 	lw	%ra, [%sp + 2]
"10010011110000010000000000000001",	-- 9663: 	lf	%f1, [%sp + 1]
"11101100001000000000000000000000",	-- 9664: 	divf	%f0, %f1, %f0
"01001111111000000000000000000000",	-- 9665: 	jr	%ra
	-- adjust_position.3000:
"11101000000000000000000000000000",	-- 9666: 	mulf	%f0, %f0, %f0
"00010100000000101100110011001101",	-- 9667: 	llif	%f2, 0.100000
"00010000000000100011110111001100",	-- 9668: 	lhif	%f2, 0.100000
"11100000000000100000000000000000",	-- 9669: 	addf	%f0, %f0, %f2
"10110000001111100000000000000000",	-- 9670: 	sf	%f1, [%sp + 0]
"00111111111111100000000000000001",	-- 9671: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 9672: 	addi	%sp, %sp, 2
"01011000000000000010101000101110",	-- 9673: 	jal	yj_sqrt
"10101011110111100000000000000010",	-- 9674: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 9675: 	lw	%ra, [%sp + 1]
"00010100000000010000000000000000",	-- 9676: 	llif	%f1, 1.000000
"00010000000000010011111110000000",	-- 9677: 	lhif	%f1, 1.000000
"11101100001000000000100000000000",	-- 9678: 	divf	%f1, %f1, %f0
"10110000000111100000000000000001",	-- 9679: 	sf	%f0, [%sp + 1]
"00001100001000000000000000000000",	-- 9680: 	movf	%f0, %f1
"00111111111111100000000000000010",	-- 9681: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9682: 	addi	%sp, %sp, 3
"01011000000000000000010010011100",	-- 9683: 	jal	atan.2520
"10101011110111100000000000000011",	-- 9684: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9685: 	lw	%ra, [%sp + 2]
"10010011110000010000000000000000",	-- 9686: 	lf	%f1, [%sp + 0]
"11101000000000010000000000000000",	-- 9687: 	mulf	%f0, %f0, %f1
"00111111111111100000000000000010",	-- 9688: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9689: 	addi	%sp, %sp, 3
"01011000000000000010010110110001",	-- 9690: 	jal	tan.2998
"10101011110111100000000000000011",	-- 9691: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9692: 	lw	%ra, [%sp + 2]
"10010011110000010000000000000001",	-- 9693: 	lf	%f1, [%sp + 1]
"11101000000000010000000000000000",	-- 9694: 	mulf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 9695: 	jr	%ra
	-- calc_dirvec.3003:
"00111011011001000000000000000001",	-- 9696: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000101",	-- 9697: 	lli	%r5, 5
"00110000101000010000000011011111",	-- 9698: 	bgt	%r5, %r1, bgt_else.9266
"00111100011111100000000000000000",	-- 9699: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 9700: 	sw	%r2, [%sp + 1]
"00111100100111100000000000000010",	-- 9701: 	sw	%r4, [%sp + 2]
"10110000000111100000000000000011",	-- 9702: 	sf	%f0, [%sp + 3]
"10110000001111100000000000000100",	-- 9703: 	sf	%f1, [%sp + 4]
"00111111111111100000000000000101",	-- 9704: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 9705: 	addi	%sp, %sp, 6
"01011000000000000000010011101111",	-- 9706: 	jal	fsqr.2530
"10101011110111100000000000000110",	-- 9707: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 9708: 	lw	%ra, [%sp + 5]
"10010011110000010000000000000100",	-- 9709: 	lf	%f1, [%sp + 4]
"10110000000111100000000000000101",	-- 9710: 	sf	%f0, [%sp + 5]
"00001100001000000000000000000000",	-- 9711: 	movf	%f0, %f1
"00111111111111100000000000000110",	-- 9712: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 9713: 	addi	%sp, %sp, 7
"01011000000000000000010011101111",	-- 9714: 	jal	fsqr.2530
"10101011110111100000000000000111",	-- 9715: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 9716: 	lw	%ra, [%sp + 6]
"10010011110000010000000000000101",	-- 9717: 	lf	%f1, [%sp + 5]
"11100000001000000000000000000000",	-- 9718: 	addf	%f0, %f1, %f0
"00010100000000010000000000000000",	-- 9719: 	llif	%f1, 1.000000
"00010000000000010011111110000000",	-- 9720: 	lhif	%f1, 1.000000
"11100000000000010000000000000000",	-- 9721: 	addf	%f0, %f0, %f1
"00111111111111100000000000000110",	-- 9722: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 9723: 	addi	%sp, %sp, 7
"01011000000000000010101000101110",	-- 9724: 	jal	yj_sqrt
"10101011110111100000000000000111",	-- 9725: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 9726: 	lw	%ra, [%sp + 6]
"10010011110000010000000000000011",	-- 9727: 	lf	%f1, [%sp + 3]
"11101100001000000000100000000000",	-- 9728: 	divf	%f1, %f1, %f0
"10010011110000100000000000000100",	-- 9729: 	lf	%f2, [%sp + 4]
"11101100010000000001000000000000",	-- 9730: 	divf	%f2, %f2, %f0
"00010100000000110000000000000000",	-- 9731: 	llif	%f3, 1.000000
"00010000000000110011111110000000",	-- 9732: 	lhif	%f3, 1.000000
"11101100011000000000000000000000",	-- 9733: 	divf	%f0, %f3, %f0
"00111011110000010000000000000001",	-- 9734: 	lw	%r1, [%sp + 1]
"00111011110000100000000000000010",	-- 9735: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 9736: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 9737: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000000000",	-- 9738: 	lw	%r2, [%sp + 0]
"10000100001000100001100000000000",	-- 9739: 	add	%r3, %r1, %r2
"00111000011000110000000000000000",	-- 9740: 	lw	%r3, [%r3 + 0]
"00111100001111100000000000000110",	-- 9741: 	sw	%r1, [%sp + 6]
"10110000000111100000000000000111",	-- 9742: 	sf	%f0, [%sp + 7]
"10110000010111100000000000001000",	-- 9743: 	sf	%f2, [%sp + 8]
"10110000001111100000000000001001",	-- 9744: 	sf	%f1, [%sp + 9]
"10000100000000110000100000000000",	-- 9745: 	add	%r1, %r0, %r3
"00111111111111100000000000001010",	-- 9746: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 9747: 	addi	%sp, %sp, 11
"01011000000000000000011010111010",	-- 9748: 	jal	d_vec.2683
"10101011110111100000000000001011",	-- 9749: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 9750: 	lw	%ra, [%sp + 10]
"10010011110000000000000000001001",	-- 9751: 	lf	%f0, [%sp + 9]
"10010011110000010000000000001000",	-- 9752: 	lf	%f1, [%sp + 8]
"10010011110000100000000000000111",	-- 9753: 	lf	%f2, [%sp + 7]
"00111111111111100000000000001010",	-- 9754: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 9755: 	addi	%sp, %sp, 11
"01011000000000000000010100100100",	-- 9756: 	jal	vecset.2576
"10101011110111100000000000001011",	-- 9757: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 9758: 	lw	%ra, [%sp + 10]
"11001100000000010000000000101000",	-- 9759: 	lli	%r1, 40
"00111011110000100000000000000000",	-- 9760: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 9761: 	add	%r1, %r2, %r1
"00111011110000110000000000000110",	-- 9762: 	lw	%r3, [%sp + 6]
"10000100011000010000100000000000",	-- 9763: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 9764: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001010",	-- 9765: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 9766: 	addi	%sp, %sp, 11
"01011000000000000000011010111010",	-- 9767: 	jal	d_vec.2683
"10101011110111100000000000001011",	-- 9768: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 9769: 	lw	%ra, [%sp + 10]
"10010011110000000000000000001000",	-- 9770: 	lf	%f0, [%sp + 8]
"00111100001111100000000000001010",	-- 9771: 	sw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 9772: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 9773: 	addi	%sp, %sp, 12
"01011000000000000010101001001111",	-- 9774: 	jal	yj_fneg
"10101011110111100000000000001100",	-- 9775: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9776: 	lw	%ra, [%sp + 11]
"00001100000000100000000000000000",	-- 9777: 	movf	%f2, %f0
"10010011110000000000000000001001",	-- 9778: 	lf	%f0, [%sp + 9]
"10010011110000010000000000000111",	-- 9779: 	lf	%f1, [%sp + 7]
"00111011110000010000000000001010",	-- 9780: 	lw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 9781: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 9782: 	addi	%sp, %sp, 12
"01011000000000000000010100100100",	-- 9783: 	jal	vecset.2576
"10101011110111100000000000001100",	-- 9784: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9785: 	lw	%ra, [%sp + 11]
"11001100000000010000000001010000",	-- 9786: 	lli	%r1, 80
"00111011110000100000000000000000",	-- 9787: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 9788: 	add	%r1, %r2, %r1
"00111011110000110000000000000110",	-- 9789: 	lw	%r3, [%sp + 6]
"10000100011000010000100000000000",	-- 9790: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 9791: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001011",	-- 9792: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 9793: 	addi	%sp, %sp, 12
"01011000000000000000011010111010",	-- 9794: 	jal	d_vec.2683
"10101011110111100000000000001100",	-- 9795: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9796: 	lw	%ra, [%sp + 11]
"10010011110000000000000000001001",	-- 9797: 	lf	%f0, [%sp + 9]
"00111100001111100000000000001011",	-- 9798: 	sw	%r1, [%sp + 11]
"00111111111111100000000000001100",	-- 9799: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 9800: 	addi	%sp, %sp, 13
"01011000000000000010101001001111",	-- 9801: 	jal	yj_fneg
"10101011110111100000000000001101",	-- 9802: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 9803: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001000",	-- 9804: 	lf	%f1, [%sp + 8]
"10110000000111100000000000001100",	-- 9805: 	sf	%f0, [%sp + 12]
"00001100001000000000000000000000",	-- 9806: 	movf	%f0, %f1
"00111111111111100000000000001101",	-- 9807: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 9808: 	addi	%sp, %sp, 14
"01011000000000000010101001001111",	-- 9809: 	jal	yj_fneg
"10101011110111100000000000001110",	-- 9810: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 9811: 	lw	%ra, [%sp + 13]
"00001100000000100000000000000000",	-- 9812: 	movf	%f2, %f0
"10010011110000000000000000000111",	-- 9813: 	lf	%f0, [%sp + 7]
"10010011110000010000000000001100",	-- 9814: 	lf	%f1, [%sp + 12]
"00111011110000010000000000001011",	-- 9815: 	lw	%r1, [%sp + 11]
"00111111111111100000000000001101",	-- 9816: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 9817: 	addi	%sp, %sp, 14
"01011000000000000000010100100100",	-- 9818: 	jal	vecset.2576
"10101011110111100000000000001110",	-- 9819: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 9820: 	lw	%ra, [%sp + 13]
"11001100000000010000000000000001",	-- 9821: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 9822: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 9823: 	add	%r1, %r2, %r1
"00111011110000110000000000000110",	-- 9824: 	lw	%r3, [%sp + 6]
"10000100011000010000100000000000",	-- 9825: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 9826: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001101",	-- 9827: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 9828: 	addi	%sp, %sp, 14
"01011000000000000000011010111010",	-- 9829: 	jal	d_vec.2683
"10101011110111100000000000001110",	-- 9830: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 9831: 	lw	%ra, [%sp + 13]
"10010011110000000000000000001001",	-- 9832: 	lf	%f0, [%sp + 9]
"00111100001111100000000000001101",	-- 9833: 	sw	%r1, [%sp + 13]
"00111111111111100000000000001110",	-- 9834: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 9835: 	addi	%sp, %sp, 15
"01011000000000000010101001001111",	-- 9836: 	jal	yj_fneg
"10101011110111100000000000001111",	-- 9837: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 9838: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001000",	-- 9839: 	lf	%f1, [%sp + 8]
"10110000000111100000000000001110",	-- 9840: 	sf	%f0, [%sp + 14]
"00001100001000000000000000000000",	-- 9841: 	movf	%f0, %f1
"00111111111111100000000000001111",	-- 9842: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9843: 	addi	%sp, %sp, 16
"01011000000000000010101001001111",	-- 9844: 	jal	yj_fneg
"10101011110111100000000000010000",	-- 9845: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9846: 	lw	%ra, [%sp + 15]
"10010011110000010000000000000111",	-- 9847: 	lf	%f1, [%sp + 7]
"10110000000111100000000000001111",	-- 9848: 	sf	%f0, [%sp + 15]
"00001100001000000000000000000000",	-- 9849: 	movf	%f0, %f1
"00111111111111100000000000010000",	-- 9850: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 9851: 	addi	%sp, %sp, 17
"01011000000000000010101001001111",	-- 9852: 	jal	yj_fneg
"10101011110111100000000000010001",	-- 9853: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 9854: 	lw	%ra, [%sp + 16]
"00001100000000100000000000000000",	-- 9855: 	movf	%f2, %f0
"10010011110000000000000000001110",	-- 9856: 	lf	%f0, [%sp + 14]
"10010011110000010000000000001111",	-- 9857: 	lf	%f1, [%sp + 15]
"00111011110000010000000000001101",	-- 9858: 	lw	%r1, [%sp + 13]
"00111111111111100000000000010000",	-- 9859: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 9860: 	addi	%sp, %sp, 17
"01011000000000000000010100100100",	-- 9861: 	jal	vecset.2576
"10101011110111100000000000010001",	-- 9862: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 9863: 	lw	%ra, [%sp + 16]
"11001100000000010000000000101001",	-- 9864: 	lli	%r1, 41
"00111011110000100000000000000000",	-- 9865: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 9866: 	add	%r1, %r2, %r1
"00111011110000110000000000000110",	-- 9867: 	lw	%r3, [%sp + 6]
"10000100011000010000100000000000",	-- 9868: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 9869: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000010000",	-- 9870: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 9871: 	addi	%sp, %sp, 17
"01011000000000000000011010111010",	-- 9872: 	jal	d_vec.2683
"10101011110111100000000000010001",	-- 9873: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 9874: 	lw	%ra, [%sp + 16]
"10010011110000000000000000001001",	-- 9875: 	lf	%f0, [%sp + 9]
"00111100001111100000000000010000",	-- 9876: 	sw	%r1, [%sp + 16]
"00111111111111100000000000010001",	-- 9877: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 9878: 	addi	%sp, %sp, 18
"01011000000000000010101001001111",	-- 9879: 	jal	yj_fneg
"10101011110111100000000000010010",	-- 9880: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 9881: 	lw	%ra, [%sp + 17]
"10010011110000010000000000000111",	-- 9882: 	lf	%f1, [%sp + 7]
"10110000000111100000000000010001",	-- 9883: 	sf	%f0, [%sp + 17]
"00001100001000000000000000000000",	-- 9884: 	movf	%f0, %f1
"00111111111111100000000000010010",	-- 9885: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 9886: 	addi	%sp, %sp, 19
"01011000000000000010101001001111",	-- 9887: 	jal	yj_fneg
"10101011110111100000000000010011",	-- 9888: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 9889: 	lw	%ra, [%sp + 18]
"00001100000000010000000000000000",	-- 9890: 	movf	%f1, %f0
"10010011110000000000000000010001",	-- 9891: 	lf	%f0, [%sp + 17]
"10010011110000100000000000001000",	-- 9892: 	lf	%f2, [%sp + 8]
"00111011110000010000000000010000",	-- 9893: 	lw	%r1, [%sp + 16]
"00111111111111100000000000010010",	-- 9894: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 9895: 	addi	%sp, %sp, 19
"01011000000000000000010100100100",	-- 9896: 	jal	vecset.2576
"10101011110111100000000000010011",	-- 9897: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 9898: 	lw	%ra, [%sp + 18]
"11001100000000010000000001010001",	-- 9899: 	lli	%r1, 81
"00111011110000100000000000000000",	-- 9900: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 9901: 	add	%r1, %r2, %r1
"00111011110000100000000000000110",	-- 9902: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 9903: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 9904: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000010010",	-- 9905: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 9906: 	addi	%sp, %sp, 19
"01011000000000000000011010111010",	-- 9907: 	jal	d_vec.2683
"10101011110111100000000000010011",	-- 9908: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 9909: 	lw	%ra, [%sp + 18]
"10010011110000000000000000000111",	-- 9910: 	lf	%f0, [%sp + 7]
"00111100001111100000000000010010",	-- 9911: 	sw	%r1, [%sp + 18]
"00111111111111100000000000010011",	-- 9912: 	sw	%ra, [%sp + 19]
"10100111110111100000000000010100",	-- 9913: 	addi	%sp, %sp, 20
"01011000000000000010101001001111",	-- 9914: 	jal	yj_fneg
"10101011110111100000000000010100",	-- 9915: 	subi	%sp, %sp, 20
"00111011110111110000000000010011",	-- 9916: 	lw	%ra, [%sp + 19]
"10010011110000010000000000001001",	-- 9917: 	lf	%f1, [%sp + 9]
"10010011110000100000000000001000",	-- 9918: 	lf	%f2, [%sp + 8]
"00111011110000010000000000010010",	-- 9919: 	lw	%r1, [%sp + 18]
"01010100000000000000010100100100",	-- 9920: 	j	vecset.2576
	-- bgt_else.9266:
"10110000010111100000000000010011",	-- 9921: 	sf	%f2, [%sp + 19]
"00111100011111100000000000000000",	-- 9922: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 9923: 	sw	%r2, [%sp + 1]
"00111111011111100000000000010100",	-- 9924: 	sw	%r27, [%sp + 20]
"10110000011111100000000000010101",	-- 9925: 	sf	%f3, [%sp + 21]
"00111100001111100000000000010110",	-- 9926: 	sw	%r1, [%sp + 22]
"00001100001000000000000000000000",	-- 9927: 	movf	%f0, %f1
"00001100010000010000000000000000",	-- 9928: 	movf	%f1, %f2
"00111111111111100000000000010111",	-- 9929: 	sw	%ra, [%sp + 23]
"10100111110111100000000000011000",	-- 9930: 	addi	%sp, %sp, 24
"01011000000000000010010111000010",	-- 9931: 	jal	adjust_position.3000
"10101011110111100000000000011000",	-- 9932: 	subi	%sp, %sp, 24
"00111011110111110000000000010111",	-- 9933: 	lw	%ra, [%sp + 23]
"11001100000000010000000000000001",	-- 9934: 	lli	%r1, 1
"00111011110000100000000000010110",	-- 9935: 	lw	%r2, [%sp + 22]
"10000100010000010000100000000000",	-- 9936: 	add	%r1, %r2, %r1
"10010011110000010000000000010101",	-- 9937: 	lf	%f1, [%sp + 21]
"10110000000111100000000000010111",	-- 9938: 	sf	%f0, [%sp + 23]
"00111100001111100000000000011000",	-- 9939: 	sw	%r1, [%sp + 24]
"00111111111111100000000000011001",	-- 9940: 	sw	%ra, [%sp + 25]
"10100111110111100000000000011010",	-- 9941: 	addi	%sp, %sp, 26
"01011000000000000010010111000010",	-- 9942: 	jal	adjust_position.3000
"10101011110111100000000000011010",	-- 9943: 	subi	%sp, %sp, 26
"00111011110111110000000000011001",	-- 9944: 	lw	%ra, [%sp + 25]
"00001100000000010000000000000000",	-- 9945: 	movf	%f1, %f0
"10010011110000000000000000010111",	-- 9946: 	lf	%f0, [%sp + 23]
"10010011110000100000000000010011",	-- 9947: 	lf	%f2, [%sp + 19]
"10010011110000110000000000010101",	-- 9948: 	lf	%f3, [%sp + 21]
"00111011110000010000000000011000",	-- 9949: 	lw	%r1, [%sp + 24]
"00111011110000100000000000000001",	-- 9950: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 9951: 	lw	%r3, [%sp + 0]
"00111011110110110000000000010100",	-- 9952: 	lw	%r27, [%sp + 20]
"00111011011110100000000000000000",	-- 9953: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 9954: 	jr	%r26
	-- calc_dirvecs.3011:
"00111011011001000000000000000001",	-- 9955: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 9956: 	lli	%r5, 0
"00110000101000010000000001010011",	-- 9957: 	bgt	%r5, %r1, bgt_else.9267
"00111111011111100000000000000000",	-- 9958: 	sw	%r27, [%sp + 0]
"00111100001111100000000000000001",	-- 9959: 	sw	%r1, [%sp + 1]
"10110000000111100000000000000010",	-- 9960: 	sf	%f0, [%sp + 2]
"00111100011111100000000000000011",	-- 9961: 	sw	%r3, [%sp + 3]
"00111100010111100000000000000100",	-- 9962: 	sw	%r2, [%sp + 4]
"00111100100111100000000000000101",	-- 9963: 	sw	%r4, [%sp + 5]
"00111111111111100000000000000110",	-- 9964: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 9965: 	addi	%sp, %sp, 7
"01011000000000000010101000101010",	-- 9966: 	jal	yj_float_of_int
"10101011110111100000000000000111",	-- 9967: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 9968: 	lw	%ra, [%sp + 6]
"00010100000000011100110011001101",	-- 9969: 	llif	%f1, 0.200000
"00010000000000010011111001001100",	-- 9970: 	lhif	%f1, 0.200000
"11101000000000010000000000000000",	-- 9971: 	mulf	%f0, %f0, %f1
"00010100000000010110011001100110",	-- 9972: 	llif	%f1, 0.900000
"00010000000000010011111101100110",	-- 9973: 	lhif	%f1, 0.900000
"11100100000000010001000000000000",	-- 9974: 	subf	%f2, %f0, %f1
"11001100000000010000000000000000",	-- 9975: 	lli	%r1, 0
"00010100000000000000000000000000",	-- 9976: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9977: 	lhif	%f0, 0.000000
"00010100000000010000000000000000",	-- 9978: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 9979: 	lhif	%f1, 0.000000
"10010011110000110000000000000010",	-- 9980: 	lf	%f3, [%sp + 2]
"00111011110000100000000000000100",	-- 9981: 	lw	%r2, [%sp + 4]
"00111011110000110000000000000011",	-- 9982: 	lw	%r3, [%sp + 3]
"00111011110110110000000000000101",	-- 9983: 	lw	%r27, [%sp + 5]
"00111111111111100000000000000110",	-- 9984: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 9985: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 9986: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 9987: 	jalr	%r26
"10101011110111100000000000000111",	-- 9988: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 9989: 	lw	%ra, [%sp + 6]
"00111011110000010000000000000001",	-- 9990: 	lw	%r1, [%sp + 1]
"00111111111111100000000000000110",	-- 9991: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 9992: 	addi	%sp, %sp, 7
"01011000000000000010101000101010",	-- 9993: 	jal	yj_float_of_int
"10101011110111100000000000000111",	-- 9994: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 9995: 	lw	%ra, [%sp + 6]
"00010100000000011100110011001101",	-- 9996: 	llif	%f1, 0.200000
"00010000000000010011111001001100",	-- 9997: 	lhif	%f1, 0.200000
"11101000000000010000000000000000",	-- 9998: 	mulf	%f0, %f0, %f1
"00010100000000011100110011001101",	-- 9999: 	llif	%f1, 0.100000
"00010000000000010011110111001100",	-- 10000: 	lhif	%f1, 0.100000
"11100000000000010001000000000000",	-- 10001: 	addf	%f2, %f0, %f1
"11001100000000010000000000000000",	-- 10002: 	lli	%r1, 0
"00010100000000000000000000000000",	-- 10003: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 10004: 	lhif	%f0, 0.000000
"00010100000000010000000000000000",	-- 10005: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 10006: 	lhif	%f1, 0.000000
"11001100000000100000000000000010",	-- 10007: 	lli	%r2, 2
"00111011110000110000000000000011",	-- 10008: 	lw	%r3, [%sp + 3]
"10000100011000100001000000000000",	-- 10009: 	add	%r2, %r3, %r2
"10010011110000110000000000000010",	-- 10010: 	lf	%f3, [%sp + 2]
"00111011110001000000000000000100",	-- 10011: 	lw	%r4, [%sp + 4]
"00111011110110110000000000000101",	-- 10012: 	lw	%r27, [%sp + 5]
"10000100000000100001100000000000",	-- 10013: 	add	%r3, %r0, %r2
"10000100000001000001000000000000",	-- 10014: 	add	%r2, %r0, %r4
"00111111111111100000000000000110",	-- 10015: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 10016: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 10017: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 10018: 	jalr	%r26
"10101011110111100000000000000111",	-- 10019: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 10020: 	lw	%ra, [%sp + 6]
"11001100000000010000000000000001",	-- 10021: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 10022: 	lw	%r2, [%sp + 1]
"10001000010000010000100000000000",	-- 10023: 	sub	%r1, %r2, %r1
"11001100000000100000000000000001",	-- 10024: 	lli	%r2, 1
"00111011110000110000000000000100",	-- 10025: 	lw	%r3, [%sp + 4]
"00111100001111100000000000000110",	-- 10026: 	sw	%r1, [%sp + 6]
"10000100000000110000100000000000",	-- 10027: 	add	%r1, %r0, %r3
"00111111111111100000000000000111",	-- 10028: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 10029: 	addi	%sp, %sp, 8
"01011000000000000000010100011101",	-- 10030: 	jal	add_mod5.2573
"10101011110111100000000000001000",	-- 10031: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 10032: 	lw	%ra, [%sp + 7]
"10000100000000010001000000000000",	-- 10033: 	add	%r2, %r0, %r1
"10010011110000000000000000000010",	-- 10034: 	lf	%f0, [%sp + 2]
"00111011110000010000000000000110",	-- 10035: 	lw	%r1, [%sp + 6]
"00111011110000110000000000000011",	-- 10036: 	lw	%r3, [%sp + 3]
"00111011110110110000000000000000",	-- 10037: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10038: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10039: 	jr	%r26
	-- bgt_else.9267:
"01001111111000000000000000000000",	-- 10040: 	jr	%ra
	-- calc_dirvec_rows.3016:
"00111011011001000000000000000001",	-- 10041: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 10042: 	lli	%r5, 0
"00110000101000010000000000101111",	-- 10043: 	bgt	%r5, %r1, bgt_else.9269
"00111111011111100000000000000000",	-- 10044: 	sw	%r27, [%sp + 0]
"00111100001111100000000000000001",	-- 10045: 	sw	%r1, [%sp + 1]
"00111100011111100000000000000010",	-- 10046: 	sw	%r3, [%sp + 2]
"00111100010111100000000000000011",	-- 10047: 	sw	%r2, [%sp + 3]
"00111100100111100000000000000100",	-- 10048: 	sw	%r4, [%sp + 4]
"00111111111111100000000000000101",	-- 10049: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 10050: 	addi	%sp, %sp, 6
"01011000000000000010101000101010",	-- 10051: 	jal	yj_float_of_int
"10101011110111100000000000000110",	-- 10052: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 10053: 	lw	%ra, [%sp + 5]
"00010100000000011100110011001101",	-- 10054: 	llif	%f1, 0.200000
"00010000000000010011111001001100",	-- 10055: 	lhif	%f1, 0.200000
"11101000000000010000000000000000",	-- 10056: 	mulf	%f0, %f0, %f1
"00010100000000010110011001100110",	-- 10057: 	llif	%f1, 0.900000
"00010000000000010011111101100110",	-- 10058: 	lhif	%f1, 0.900000
"11100100000000010000000000000000",	-- 10059: 	subf	%f0, %f0, %f1
"11001100000000010000000000000100",	-- 10060: 	lli	%r1, 4
"00111011110000100000000000000011",	-- 10061: 	lw	%r2, [%sp + 3]
"00111011110000110000000000000010",	-- 10062: 	lw	%r3, [%sp + 2]
"00111011110110110000000000000100",	-- 10063: 	lw	%r27, [%sp + 4]
"00111111111111100000000000000101",	-- 10064: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 10065: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 10066: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 10067: 	jalr	%r26
"10101011110111100000000000000110",	-- 10068: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 10069: 	lw	%ra, [%sp + 5]
"11001100000000010000000000000001",	-- 10070: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 10071: 	lw	%r2, [%sp + 1]
"10001000010000010000100000000000",	-- 10072: 	sub	%r1, %r2, %r1
"11001100000000100000000000000010",	-- 10073: 	lli	%r2, 2
"00111011110000110000000000000011",	-- 10074: 	lw	%r3, [%sp + 3]
"00111100001111100000000000000101",	-- 10075: 	sw	%r1, [%sp + 5]
"10000100000000110000100000000000",	-- 10076: 	add	%r1, %r0, %r3
"00111111111111100000000000000110",	-- 10077: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 10078: 	addi	%sp, %sp, 7
"01011000000000000000010100011101",	-- 10079: 	jal	add_mod5.2573
"10101011110111100000000000000111",	-- 10080: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 10081: 	lw	%ra, [%sp + 6]
"10000100000000010001000000000000",	-- 10082: 	add	%r2, %r0, %r1
"11001100000000010000000000000100",	-- 10083: 	lli	%r1, 4
"00111011110000110000000000000010",	-- 10084: 	lw	%r3, [%sp + 2]
"10000100011000010001100000000000",	-- 10085: 	add	%r3, %r3, %r1
"00111011110000010000000000000101",	-- 10086: 	lw	%r1, [%sp + 5]
"00111011110110110000000000000000",	-- 10087: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10088: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10089: 	jr	%r26
	-- bgt_else.9269:
"01001111111000000000000000000000",	-- 10090: 	jr	%ra
	-- create_dirvec.3020:
"00111011011000010000000000000001",	-- 10091: 	lw	%r1, [%r27 + 1]
"11001100000000100000000000000011",	-- 10092: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 10093: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 10094: 	lhif	%f0, 0.000000
"00111100001111100000000000000000",	-- 10095: 	sw	%r1, [%sp + 0]
"10000100000000100000100000000000",	-- 10096: 	add	%r1, %r0, %r2
"00111111111111100000000000000001",	-- 10097: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 10098: 	addi	%sp, %sp, 2
"01011000000000000010101000100010",	-- 10099: 	jal	yj_create_float_array
"10101011110111100000000000000010",	-- 10100: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 10101: 	lw	%ra, [%sp + 1]
"10000100000000010001000000000000",	-- 10102: 	add	%r2, %r0, %r1
"11001100000000010000000000000000",	-- 10103: 	lli	%r1, 0
"00111011110000110000000000000000",	-- 10104: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 10105: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 10106: 	lw	%r1, [%r1 + 0]
"00111100010111100000000000000001",	-- 10107: 	sw	%r2, [%sp + 1]
"00111111111111100000000000000010",	-- 10108: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 10109: 	addi	%sp, %sp, 3
"01011000000000000010101000011010",	-- 10110: 	jal	yj_create_array
"10101011110111100000000000000011",	-- 10111: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 10112: 	lw	%ra, [%sp + 2]
"10000100000111010001000000000000",	-- 10113: 	add	%r2, %r0, %hp
"10100111101111010000000000000010",	-- 10114: 	addi	%hp, %hp, 2
"00111100001000100000000000000001",	-- 10115: 	sw	%r1, [%r2 + 1]
"00111011110000010000000000000001",	-- 10116: 	lw	%r1, [%sp + 1]
"00111100001000100000000000000000",	-- 10117: 	sw	%r1, [%r2 + 0]
"10000100000000100000100000000000",	-- 10118: 	add	%r1, %r0, %r2
"01001111111000000000000000000000",	-- 10119: 	jr	%ra
	-- create_dirvec_elements.3022:
"00111011011000110000000000000001",	-- 10120: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 10121: 	lli	%r4, 0
"00110000100000100000000000010101",	-- 10122: 	bgt	%r4, %r2, bgt_else.9271
"00111111011111100000000000000000",	-- 10123: 	sw	%r27, [%sp + 0]
"00111100010111100000000000000001",	-- 10124: 	sw	%r2, [%sp + 1]
"00111100001111100000000000000010",	-- 10125: 	sw	%r1, [%sp + 2]
"10000100000000111101100000000000",	-- 10126: 	add	%r27, %r0, %r3
"00111111111111100000000000000011",	-- 10127: 	sw	%ra, [%sp + 3]
"00111011011110100000000000000000",	-- 10128: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000100",	-- 10129: 	addi	%sp, %sp, 4
"01010011010000000000000000000000",	-- 10130: 	jalr	%r26
"10101011110111100000000000000100",	-- 10131: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 10132: 	lw	%ra, [%sp + 3]
"00111011110000100000000000000001",	-- 10133: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000010",	-- 10134: 	lw	%r3, [%sp + 2]
"10000100011000100010000000000000",	-- 10135: 	add	%r4, %r3, %r2
"00111100001001000000000000000000",	-- 10136: 	sw	%r1, [%r4 + 0]
"11001100000000010000000000000001",	-- 10137: 	lli	%r1, 1
"10001000010000010001000000000000",	-- 10138: 	sub	%r2, %r2, %r1
"00111011110110110000000000000000",	-- 10139: 	lw	%r27, [%sp + 0]
"10000100000000110000100000000000",	-- 10140: 	add	%r1, %r0, %r3
"00111011011110100000000000000000",	-- 10141: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10142: 	jr	%r26
	-- bgt_else.9271:
"01001111111000000000000000000000",	-- 10143: 	jr	%ra
	-- create_dirvecs.3025:
"00111011011000100000000000000011",	-- 10144: 	lw	%r2, [%r27 + 3]
"00111011011000110000000000000010",	-- 10145: 	lw	%r3, [%r27 + 2]
"00111011011001000000000000000001",	-- 10146: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 10147: 	lli	%r5, 0
"00110000101000010000000000101010",	-- 10148: 	bgt	%r5, %r1, bgt_else.9273
"11001100000001010000000001111000",	-- 10149: 	lli	%r5, 120
"00111111011111100000000000000000",	-- 10150: 	sw	%r27, [%sp + 0]
"00111100011111100000000000000001",	-- 10151: 	sw	%r3, [%sp + 1]
"00111100001111100000000000000010",	-- 10152: 	sw	%r1, [%sp + 2]
"00111100010111100000000000000011",	-- 10153: 	sw	%r2, [%sp + 3]
"00111100101111100000000000000100",	-- 10154: 	sw	%r5, [%sp + 4]
"10000100000001001101100000000000",	-- 10155: 	add	%r27, %r0, %r4
"00111111111111100000000000000101",	-- 10156: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 10157: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 10158: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 10159: 	jalr	%r26
"10101011110111100000000000000110",	-- 10160: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 10161: 	lw	%ra, [%sp + 5]
"10000100000000010001000000000000",	-- 10162: 	add	%r2, %r0, %r1
"00111011110000010000000000000100",	-- 10163: 	lw	%r1, [%sp + 4]
"00111111111111100000000000000101",	-- 10164: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 10165: 	addi	%sp, %sp, 6
"01011000000000000010101000011010",	-- 10166: 	jal	yj_create_array
"10101011110111100000000000000110",	-- 10167: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 10168: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000010",	-- 10169: 	lw	%r2, [%sp + 2]
"00111011110000110000000000000011",	-- 10170: 	lw	%r3, [%sp + 3]
"10000100011000100010000000000000",	-- 10171: 	add	%r4, %r3, %r2
"00111100001001000000000000000000",	-- 10172: 	sw	%r1, [%r4 + 0]
"10000100011000100000100000000000",	-- 10173: 	add	%r1, %r3, %r2
"00111000001000010000000000000000",	-- 10174: 	lw	%r1, [%r1 + 0]
"11001100000000110000000001110110",	-- 10175: 	lli	%r3, 118
"00111011110110110000000000000001",	-- 10176: 	lw	%r27, [%sp + 1]
"10000100000000110001000000000000",	-- 10177: 	add	%r2, %r0, %r3
"00111111111111100000000000000101",	-- 10178: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 10179: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 10180: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 10181: 	jalr	%r26
"10101011110111100000000000000110",	-- 10182: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 10183: 	lw	%ra, [%sp + 5]
"11001100000000010000000000000001",	-- 10184: 	lli	%r1, 1
"00111011110000100000000000000010",	-- 10185: 	lw	%r2, [%sp + 2]
"10001000010000010000100000000000",	-- 10186: 	sub	%r1, %r2, %r1
"00111011110110110000000000000000",	-- 10187: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10188: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10189: 	jr	%r26
	-- bgt_else.9273:
"01001111111000000000000000000000",	-- 10190: 	jr	%ra
	-- init_dirvec_constants.3027:
"00111011011000110000000000000001",	-- 10191: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 10192: 	lli	%r4, 0
"00110000100000100000000000010101",	-- 10193: 	bgt	%r4, %r2, bgt_else.9275
"10000100001000100010000000000000",	-- 10194: 	add	%r4, %r1, %r2
"00111000100001000000000000000000",	-- 10195: 	lw	%r4, [%r4 + 0]
"00111100001111100000000000000000",	-- 10196: 	sw	%r1, [%sp + 0]
"00111111011111100000000000000001",	-- 10197: 	sw	%r27, [%sp + 1]
"00111100010111100000000000000010",	-- 10198: 	sw	%r2, [%sp + 2]
"10000100000001000000100000000000",	-- 10199: 	add	%r1, %r0, %r4
"10000100000000111101100000000000",	-- 10200: 	add	%r27, %r0, %r3
"00111111111111100000000000000011",	-- 10201: 	sw	%ra, [%sp + 3]
"00111011011110100000000000000000",	-- 10202: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000100",	-- 10203: 	addi	%sp, %sp, 4
"01010011010000000000000000000000",	-- 10204: 	jalr	%r26
"10101011110111100000000000000100",	-- 10205: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 10206: 	lw	%ra, [%sp + 3]
"11001100000000010000000000000001",	-- 10207: 	lli	%r1, 1
"00111011110000100000000000000010",	-- 10208: 	lw	%r2, [%sp + 2]
"10001000010000010001000000000000",	-- 10209: 	sub	%r2, %r2, %r1
"00111011110000010000000000000000",	-- 10210: 	lw	%r1, [%sp + 0]
"00111011110110110000000000000001",	-- 10211: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 10212: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10213: 	jr	%r26
	-- bgt_else.9275:
"01001111111000000000000000000000",	-- 10214: 	jr	%ra
	-- init_vecset_constants.3030:
"00111011011000100000000000000010",	-- 10215: 	lw	%r2, [%r27 + 2]
"00111011011000110000000000000001",	-- 10216: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 10217: 	lli	%r4, 0
"00110000100000010000000000010101",	-- 10218: 	bgt	%r4, %r1, bgt_else.9277
"10000100011000010001100000000000",	-- 10219: 	add	%r3, %r3, %r1
"00111000011000110000000000000000",	-- 10220: 	lw	%r3, [%r3 + 0]
"11001100000001000000000001110111",	-- 10221: 	lli	%r4, 119
"00111111011111100000000000000000",	-- 10222: 	sw	%r27, [%sp + 0]
"00111100001111100000000000000001",	-- 10223: 	sw	%r1, [%sp + 1]
"10000100000000110000100000000000",	-- 10224: 	add	%r1, %r0, %r3
"10000100000000101101100000000000",	-- 10225: 	add	%r27, %r0, %r2
"10000100000001000001000000000000",	-- 10226: 	add	%r2, %r0, %r4
"00111111111111100000000000000010",	-- 10227: 	sw	%ra, [%sp + 2]
"00111011011110100000000000000000",	-- 10228: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000011",	-- 10229: 	addi	%sp, %sp, 3
"01010011010000000000000000000000",	-- 10230: 	jalr	%r26
"10101011110111100000000000000011",	-- 10231: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 10232: 	lw	%ra, [%sp + 2]
"11001100000000010000000000000001",	-- 10233: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 10234: 	lw	%r2, [%sp + 1]
"10001000010000010000100000000000",	-- 10235: 	sub	%r1, %r2, %r1
"00111011110110110000000000000000",	-- 10236: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10237: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10238: 	jr	%r26
	-- bgt_else.9277:
"01001111111000000000000000000000",	-- 10239: 	jr	%ra
	-- init_dirvecs.3032:
"00111011011000010000000000000011",	-- 10240: 	lw	%r1, [%r27 + 3]
"00111011011000100000000000000010",	-- 10241: 	lw	%r2, [%r27 + 2]
"00111011011000110000000000000001",	-- 10242: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000100",	-- 10243: 	lli	%r4, 4
"00111100001111100000000000000000",	-- 10244: 	sw	%r1, [%sp + 0]
"00111100011111100000000000000001",	-- 10245: 	sw	%r3, [%sp + 1]
"10000100000001000000100000000000",	-- 10246: 	add	%r1, %r0, %r4
"10000100000000101101100000000000",	-- 10247: 	add	%r27, %r0, %r2
"00111111111111100000000000000010",	-- 10248: 	sw	%ra, [%sp + 2]
"00111011011110100000000000000000",	-- 10249: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000011",	-- 10250: 	addi	%sp, %sp, 3
"01010011010000000000000000000000",	-- 10251: 	jalr	%r26
"10101011110111100000000000000011",	-- 10252: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 10253: 	lw	%ra, [%sp + 2]
"11001100000000010000000000001001",	-- 10254: 	lli	%r1, 9
"11001100000000100000000000000000",	-- 10255: 	lli	%r2, 0
"11001100000000110000000000000000",	-- 10256: 	lli	%r3, 0
"00111011110110110000000000000001",	-- 10257: 	lw	%r27, [%sp + 1]
"00111111111111100000000000000010",	-- 10258: 	sw	%ra, [%sp + 2]
"00111011011110100000000000000000",	-- 10259: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000011",	-- 10260: 	addi	%sp, %sp, 3
"01010011010000000000000000000000",	-- 10261: 	jalr	%r26
"10101011110111100000000000000011",	-- 10262: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 10263: 	lw	%ra, [%sp + 2]
"11001100000000010000000000000100",	-- 10264: 	lli	%r1, 4
"00111011110110110000000000000000",	-- 10265: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10266: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10267: 	jr	%r26
	-- add_reflection.3034:
"00111011011000110000000000000011",	-- 10268: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 10269: 	lw	%r4, [%r27 + 2]
"00111011011110110000000000000001",	-- 10270: 	lw	%r27, [%r27 + 1]
"00111100001111100000000000000000",	-- 10271: 	sw	%r1, [%sp + 0]
"00111100100111100000000000000001",	-- 10272: 	sw	%r4, [%sp + 1]
"00111100010111100000000000000010",	-- 10273: 	sw	%r2, [%sp + 2]
"10110000000111100000000000000011",	-- 10274: 	sf	%f0, [%sp + 3]
"00111100011111100000000000000100",	-- 10275: 	sw	%r3, [%sp + 4]
"10110000011111100000000000000101",	-- 10276: 	sf	%f3, [%sp + 5]
"10110000010111100000000000000110",	-- 10277: 	sf	%f2, [%sp + 6]
"10110000001111100000000000000111",	-- 10278: 	sf	%f1, [%sp + 7]
"00111111111111100000000000001000",	-- 10279: 	sw	%ra, [%sp + 8]
"00111011011110100000000000000000",	-- 10280: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001001",	-- 10281: 	addi	%sp, %sp, 9
"01010011010000000000000000000000",	-- 10282: 	jalr	%r26
"10101011110111100000000000001001",	-- 10283: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 10284: 	lw	%ra, [%sp + 8]
"00111100001111100000000000001000",	-- 10285: 	sw	%r1, [%sp + 8]
"00111111111111100000000000001001",	-- 10286: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 10287: 	addi	%sp, %sp, 10
"01011000000000000000011010111010",	-- 10288: 	jal	d_vec.2683
"10101011110111100000000000001010",	-- 10289: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 10290: 	lw	%ra, [%sp + 9]
"10010011110000000000000000000111",	-- 10291: 	lf	%f0, [%sp + 7]
"10010011110000010000000000000110",	-- 10292: 	lf	%f1, [%sp + 6]
"10010011110000100000000000000101",	-- 10293: 	lf	%f2, [%sp + 5]
"00111111111111100000000000001001",	-- 10294: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 10295: 	addi	%sp, %sp, 10
"01011000000000000000010100100100",	-- 10296: 	jal	vecset.2576
"10101011110111100000000000001010",	-- 10297: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 10298: 	lw	%ra, [%sp + 9]
"00111011110000010000000000001000",	-- 10299: 	lw	%r1, [%sp + 8]
"00111011110110110000000000000100",	-- 10300: 	lw	%r27, [%sp + 4]
"00111111111111100000000000001001",	-- 10301: 	sw	%ra, [%sp + 9]
"00111011011110100000000000000000",	-- 10302: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001010",	-- 10303: 	addi	%sp, %sp, 10
"01010011010000000000000000000000",	-- 10304: 	jalr	%r26
"10101011110111100000000000001010",	-- 10305: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 10306: 	lw	%ra, [%sp + 9]
"10000100000111010000100000000000",	-- 10307: 	add	%r1, %r0, %hp
"10100111101111010000000000000011",	-- 10308: 	addi	%hp, %hp, 3
"10010011110000000000000000000011",	-- 10309: 	lf	%f0, [%sp + 3]
"10110000000000010000000000000010",	-- 10310: 	sf	%f0, [%r1 + 2]
"00111011110000100000000000001000",	-- 10311: 	lw	%r2, [%sp + 8]
"00111100010000010000000000000001",	-- 10312: 	sw	%r2, [%r1 + 1]
"00111011110000100000000000000010",	-- 10313: 	lw	%r2, [%sp + 2]
"00111100010000010000000000000000",	-- 10314: 	sw	%r2, [%r1 + 0]
"00111011110000100000000000000000",	-- 10315: 	lw	%r2, [%sp + 0]
"00111011110000110000000000000001",	-- 10316: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 10317: 	add	%r2, %r3, %r2
"00111100001000100000000000000000",	-- 10318: 	sw	%r1, [%r2 + 0]
"01001111111000000000000000000000",	-- 10319: 	jr	%ra
	-- setup_rect_reflection.3041:
"00111011011000110000000000000011",	-- 10320: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 10321: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 10322: 	lw	%r5, [%r27 + 1]
"11001100000001100000000000000100",	-- 10323: 	lli	%r6, 4
"10001100001001100000100000000000",	-- 10324: 	mul	%r1, %r1, %r6
"11001100000001100000000000000000",	-- 10325: 	lli	%r6, 0
"10000100011001100011000000000000",	-- 10326: 	add	%r6, %r3, %r6
"00111000110001100000000000000000",	-- 10327: 	lw	%r6, [%r6 + 0]
"00010100000000000000000000000000",	-- 10328: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 10329: 	lhif	%f0, 1.000000
"00111100011111100000000000000000",	-- 10330: 	sw	%r3, [%sp + 0]
"00111100110111100000000000000001",	-- 10331: 	sw	%r6, [%sp + 1]
"00111100101111100000000000000010",	-- 10332: 	sw	%r5, [%sp + 2]
"00111100001111100000000000000011",	-- 10333: 	sw	%r1, [%sp + 3]
"00111100100111100000000000000100",	-- 10334: 	sw	%r4, [%sp + 4]
"10110000000111100000000000000101",	-- 10335: 	sf	%f0, [%sp + 5]
"10000100000000100000100000000000",	-- 10336: 	add	%r1, %r0, %r2
"00111111111111100000000000000110",	-- 10337: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 10338: 	addi	%sp, %sp, 7
"01011000000000000000011001111000",	-- 10339: 	jal	o_diffuse.2646
"10101011110111100000000000000111",	-- 10340: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 10341: 	lw	%ra, [%sp + 6]
"10010011110000010000000000000101",	-- 10342: 	lf	%f1, [%sp + 5]
"11100100001000000000000000000000",	-- 10343: 	subf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 10344: 	lli	%r1, 0
"00111011110000100000000000000100",	-- 10345: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 10346: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 10347: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000110",	-- 10348: 	sf	%f0, [%sp + 6]
"00001100001000000000000000000000",	-- 10349: 	movf	%f0, %f1
"00111111111111100000000000000111",	-- 10350: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 10351: 	addi	%sp, %sp, 8
"01011000000000000010101001001111",	-- 10352: 	jal	yj_fneg
"10101011110111100000000000001000",	-- 10353: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 10354: 	lw	%ra, [%sp + 7]
"11001100000000010000000000000001",	-- 10355: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 10356: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 10357: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 10358: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000111",	-- 10359: 	sf	%f0, [%sp + 7]
"00001100001000000000000000000000",	-- 10360: 	movf	%f0, %f1
"00111111111111100000000000001000",	-- 10361: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 10362: 	addi	%sp, %sp, 9
"01011000000000000010101001001111",	-- 10363: 	jal	yj_fneg
"10101011110111100000000000001001",	-- 10364: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 10365: 	lw	%ra, [%sp + 8]
"11001100000000010000000000000010",	-- 10366: 	lli	%r1, 2
"00111011110000100000000000000100",	-- 10367: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 10368: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 10369: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000001000",	-- 10370: 	sf	%f0, [%sp + 8]
"00001100001000000000000000000000",	-- 10371: 	movf	%f0, %f1
"00111111111111100000000000001001",	-- 10372: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 10373: 	addi	%sp, %sp, 10
"01011000000000000010101001001111",	-- 10374: 	jal	yj_fneg
"10101011110111100000000000001010",	-- 10375: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 10376: 	lw	%ra, [%sp + 9]
"00001100000000110000000000000000",	-- 10377: 	movf	%f3, %f0
"11001100000000010000000000000001",	-- 10378: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 10379: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 10380: 	add	%r1, %r2, %r1
"11001100000000110000000000000000",	-- 10381: 	lli	%r3, 0
"00111011110001000000000000000100",	-- 10382: 	lw	%r4, [%sp + 4]
"10000100100000110001100000000000",	-- 10383: 	add	%r3, %r4, %r3
"10010000011000010000000000000000",	-- 10384: 	lf	%f1, [%r3 + 0]
"10010011110000000000000000000110",	-- 10385: 	lf	%f0, [%sp + 6]
"10010011110000100000000000001000",	-- 10386: 	lf	%f2, [%sp + 8]
"00111011110000110000000000000001",	-- 10387: 	lw	%r3, [%sp + 1]
"00111011110110110000000000000010",	-- 10388: 	lw	%r27, [%sp + 2]
"10110000011111100000000000001001",	-- 10389: 	sf	%f3, [%sp + 9]
"10000100000000010001000000000000",	-- 10390: 	add	%r2, %r0, %r1
"10000100000000110000100000000000",	-- 10391: 	add	%r1, %r0, %r3
"00111111111111100000000000001010",	-- 10392: 	sw	%ra, [%sp + 10]
"00111011011110100000000000000000",	-- 10393: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001011",	-- 10394: 	addi	%sp, %sp, 11
"01010011010000000000000000000000",	-- 10395: 	jalr	%r26
"10101011110111100000000000001011",	-- 10396: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 10397: 	lw	%ra, [%sp + 10]
"11001100000000010000000000000001",	-- 10398: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 10399: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 10400: 	add	%r1, %r2, %r1
"11001100000000110000000000000010",	-- 10401: 	lli	%r3, 2
"00111011110001000000000000000011",	-- 10402: 	lw	%r4, [%sp + 3]
"10000100100000110001100000000000",	-- 10403: 	add	%r3, %r4, %r3
"11001100000001010000000000000001",	-- 10404: 	lli	%r5, 1
"00111011110001100000000000000100",	-- 10405: 	lw	%r6, [%sp + 4]
"10000100110001010010100000000000",	-- 10406: 	add	%r5, %r6, %r5
"10010000101000100000000000000000",	-- 10407: 	lf	%f2, [%r5 + 0]
"10010011110000000000000000000110",	-- 10408: 	lf	%f0, [%sp + 6]
"10010011110000010000000000000111",	-- 10409: 	lf	%f1, [%sp + 7]
"10010011110000110000000000001001",	-- 10410: 	lf	%f3, [%sp + 9]
"00111011110110110000000000000010",	-- 10411: 	lw	%r27, [%sp + 2]
"10000100000000110001000000000000",	-- 10412: 	add	%r2, %r0, %r3
"00111111111111100000000000001010",	-- 10413: 	sw	%ra, [%sp + 10]
"00111011011110100000000000000000",	-- 10414: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001011",	-- 10415: 	addi	%sp, %sp, 11
"01010011010000000000000000000000",	-- 10416: 	jalr	%r26
"10101011110111100000000000001011",	-- 10417: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 10418: 	lw	%ra, [%sp + 10]
"11001100000000010000000000000010",	-- 10419: 	lli	%r1, 2
"00111011110000100000000000000001",	-- 10420: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 10421: 	add	%r1, %r2, %r1
"11001100000000110000000000000011",	-- 10422: 	lli	%r3, 3
"00111011110001000000000000000011",	-- 10423: 	lw	%r4, [%sp + 3]
"10000100100000110001100000000000",	-- 10424: 	add	%r3, %r4, %r3
"11001100000001000000000000000010",	-- 10425: 	lli	%r4, 2
"00111011110001010000000000000100",	-- 10426: 	lw	%r5, [%sp + 4]
"10000100101001000010000000000000",	-- 10427: 	add	%r4, %r5, %r4
"10010000100000110000000000000000",	-- 10428: 	lf	%f3, [%r4 + 0]
"10010011110000000000000000000110",	-- 10429: 	lf	%f0, [%sp + 6]
"10010011110000010000000000000111",	-- 10430: 	lf	%f1, [%sp + 7]
"10010011110000100000000000001000",	-- 10431: 	lf	%f2, [%sp + 8]
"00111011110110110000000000000010",	-- 10432: 	lw	%r27, [%sp + 2]
"10000100000000110001000000000000",	-- 10433: 	add	%r2, %r0, %r3
"00111111111111100000000000001010",	-- 10434: 	sw	%ra, [%sp + 10]
"00111011011110100000000000000000",	-- 10435: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001011",	-- 10436: 	addi	%sp, %sp, 11
"01010011010000000000000000000000",	-- 10437: 	jalr	%r26
"10101011110111100000000000001011",	-- 10438: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 10439: 	lw	%ra, [%sp + 10]
"11001100000000010000000000000000",	-- 10440: 	lli	%r1, 0
"11001100000000100000000000000011",	-- 10441: 	lli	%r2, 3
"00111011110000110000000000000001",	-- 10442: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 10443: 	add	%r2, %r3, %r2
"00111011110000110000000000000000",	-- 10444: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 10445: 	add	%r1, %r3, %r1
"00111100010000010000000000000000",	-- 10446: 	sw	%r2, [%r1 + 0]
"01001111111000000000000000000000",	-- 10447: 	jr	%ra
	-- setup_surface_reflection.3044:
"00111011011000110000000000000011",	-- 10448: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 10449: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 10450: 	lw	%r5, [%r27 + 1]
"11001100000001100000000000000100",	-- 10451: 	lli	%r6, 4
"10001100001001100000100000000000",	-- 10452: 	mul	%r1, %r1, %r6
"11001100000001100000000000000001",	-- 10453: 	lli	%r6, 1
"10000100001001100000100000000000",	-- 10454: 	add	%r1, %r1, %r6
"11001100000001100000000000000000",	-- 10455: 	lli	%r6, 0
"10000100011001100011000000000000",	-- 10456: 	add	%r6, %r3, %r6
"00111000110001100000000000000000",	-- 10457: 	lw	%r6, [%r6 + 0]
"00010100000000000000000000000000",	-- 10458: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 10459: 	lhif	%f0, 1.000000
"00111100011111100000000000000000",	-- 10460: 	sw	%r3, [%sp + 0]
"00111100001111100000000000000001",	-- 10461: 	sw	%r1, [%sp + 1]
"00111100110111100000000000000010",	-- 10462: 	sw	%r6, [%sp + 2]
"00111100101111100000000000000011",	-- 10463: 	sw	%r5, [%sp + 3]
"00111100100111100000000000000100",	-- 10464: 	sw	%r4, [%sp + 4]
"00111100010111100000000000000101",	-- 10465: 	sw	%r2, [%sp + 5]
"10110000000111100000000000000110",	-- 10466: 	sf	%f0, [%sp + 6]
"10000100000000100000100000000000",	-- 10467: 	add	%r1, %r0, %r2
"00111111111111100000000000000111",	-- 10468: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 10469: 	addi	%sp, %sp, 8
"01011000000000000000011001111000",	-- 10470: 	jal	o_diffuse.2646
"10101011110111100000000000001000",	-- 10471: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 10472: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000110",	-- 10473: 	lf	%f1, [%sp + 6]
"11100100001000000000000000000000",	-- 10474: 	subf	%f0, %f1, %f0
"00111011110000010000000000000101",	-- 10475: 	lw	%r1, [%sp + 5]
"10110000000111100000000000000111",	-- 10476: 	sf	%f0, [%sp + 7]
"00111111111111100000000000001000",	-- 10477: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 10478: 	addi	%sp, %sp, 9
"01011000000000000000011001100111",	-- 10479: 	jal	o_param_abc.2638
"10101011110111100000000000001001",	-- 10480: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 10481: 	lw	%ra, [%sp + 8]
"10000100000000010001000000000000",	-- 10482: 	add	%r2, %r0, %r1
"00111011110000010000000000000100",	-- 10483: 	lw	%r1, [%sp + 4]
"00111111111111100000000000001000",	-- 10484: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 10485: 	addi	%sp, %sp, 9
"01011000000000000000010110100101",	-- 10486: 	jal	veciprod.2597
"10101011110111100000000000001001",	-- 10487: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 10488: 	lw	%ra, [%sp + 8]
"00010100000000010000000000000000",	-- 10489: 	llif	%f1, 2.000000
"00010000000000010100000000000000",	-- 10490: 	lhif	%f1, 2.000000
"00111011110000010000000000000101",	-- 10491: 	lw	%r1, [%sp + 5]
"10110000000111100000000000001000",	-- 10492: 	sf	%f0, [%sp + 8]
"10110000001111100000000000001001",	-- 10493: 	sf	%f1, [%sp + 9]
"00111111111111100000000000001010",	-- 10494: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 10495: 	addi	%sp, %sp, 11
"01011000000000000000011001011000",	-- 10496: 	jal	o_param_a.2632
"10101011110111100000000000001011",	-- 10497: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 10498: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 10499: 	lf	%f1, [%sp + 9]
"11101000001000000000000000000000",	-- 10500: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001000",	-- 10501: 	lf	%f1, [%sp + 8]
"11101000000000010000000000000000",	-- 10502: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000000",	-- 10503: 	lli	%r1, 0
"00111011110000100000000000000100",	-- 10504: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 10505: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 10506: 	lf	%f2, [%r1 + 0]
"11100100000000100000000000000000",	-- 10507: 	subf	%f0, %f0, %f2
"00010100000000100000000000000000",	-- 10508: 	llif	%f2, 2.000000
"00010000000000100100000000000000",	-- 10509: 	lhif	%f2, 2.000000
"00111011110000010000000000000101",	-- 10510: 	lw	%r1, [%sp + 5]
"10110000000111100000000000001010",	-- 10511: 	sf	%f0, [%sp + 10]
"10110000010111100000000000001011",	-- 10512: 	sf	%f2, [%sp + 11]
"00111111111111100000000000001100",	-- 10513: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 10514: 	addi	%sp, %sp, 13
"01011000000000000000011001011101",	-- 10515: 	jal	o_param_b.2634
"10101011110111100000000000001101",	-- 10516: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 10517: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001011",	-- 10518: 	lf	%f1, [%sp + 11]
"11101000001000000000000000000000",	-- 10519: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001000",	-- 10520: 	lf	%f1, [%sp + 8]
"11101000000000010000000000000000",	-- 10521: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000001",	-- 10522: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 10523: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 10524: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 10525: 	lf	%f2, [%r1 + 0]
"11100100000000100000000000000000",	-- 10526: 	subf	%f0, %f0, %f2
"00010100000000100000000000000000",	-- 10527: 	llif	%f2, 2.000000
"00010000000000100100000000000000",	-- 10528: 	lhif	%f2, 2.000000
"00111011110000010000000000000101",	-- 10529: 	lw	%r1, [%sp + 5]
"10110000000111100000000000001100",	-- 10530: 	sf	%f0, [%sp + 12]
"10110000010111100000000000001101",	-- 10531: 	sf	%f2, [%sp + 13]
"00111111111111100000000000001110",	-- 10532: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 10533: 	addi	%sp, %sp, 15
"01011000000000000000011001100010",	-- 10534: 	jal	o_param_c.2636
"10101011110111100000000000001111",	-- 10535: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 10536: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001101",	-- 10537: 	lf	%f1, [%sp + 13]
"11101000001000000000000000000000",	-- 10538: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001000",	-- 10539: 	lf	%f1, [%sp + 8]
"11101000000000010000000000000000",	-- 10540: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000010",	-- 10541: 	lli	%r1, 2
"00111011110000100000000000000100",	-- 10542: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 10543: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 10544: 	lf	%f1, [%r1 + 0]
"11100100000000010001100000000000",	-- 10545: 	subf	%f3, %f0, %f1
"10010011110000000000000000000111",	-- 10546: 	lf	%f0, [%sp + 7]
"10010011110000010000000000001010",	-- 10547: 	lf	%f1, [%sp + 10]
"10010011110000100000000000001100",	-- 10548: 	lf	%f2, [%sp + 12]
"00111011110000010000000000000010",	-- 10549: 	lw	%r1, [%sp + 2]
"00111011110000100000000000000001",	-- 10550: 	lw	%r2, [%sp + 1]
"00111011110110110000000000000011",	-- 10551: 	lw	%r27, [%sp + 3]
"00111111111111100000000000001110",	-- 10552: 	sw	%ra, [%sp + 14]
"00111011011110100000000000000000",	-- 10553: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001111",	-- 10554: 	addi	%sp, %sp, 15
"01010011010000000000000000000000",	-- 10555: 	jalr	%r26
"10101011110111100000000000001111",	-- 10556: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 10557: 	lw	%ra, [%sp + 14]
"11001100000000010000000000000000",	-- 10558: 	lli	%r1, 0
"11001100000000100000000000000001",	-- 10559: 	lli	%r2, 1
"00111011110000110000000000000010",	-- 10560: 	lw	%r3, [%sp + 2]
"10000100011000100001000000000000",	-- 10561: 	add	%r2, %r3, %r2
"00111011110000110000000000000000",	-- 10562: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 10563: 	add	%r1, %r3, %r1
"00111100010000010000000000000000",	-- 10564: 	sw	%r2, [%r1 + 0]
"01001111111000000000000000000000",	-- 10565: 	jr	%ra
	-- setup_reflections.3047:
"00111011011000100000000000000011",	-- 10566: 	lw	%r2, [%r27 + 3]
"00111011011000110000000000000010",	-- 10567: 	lw	%r3, [%r27 + 2]
"00111011011001000000000000000001",	-- 10568: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 10569: 	lli	%r5, 0
"00110000101000010000000000110101",	-- 10570: 	bgt	%r5, %r1, bgt_else.9282
"10000100100000010010000000000000",	-- 10571: 	add	%r4, %r4, %r1
"00111000100001000000000000000000",	-- 10572: 	lw	%r4, [%r4 + 0]
"00111100010111100000000000000000",	-- 10573: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 10574: 	sw	%r1, [%sp + 1]
"00111100011111100000000000000010",	-- 10575: 	sw	%r3, [%sp + 2]
"00111100100111100000000000000011",	-- 10576: 	sw	%r4, [%sp + 3]
"10000100000001000000100000000000",	-- 10577: 	add	%r1, %r0, %r4
"00111111111111100000000000000100",	-- 10578: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 10579: 	addi	%sp, %sp, 5
"01011000000000000000011001010010",	-- 10580: 	jal	o_reflectiontype.2626
"10101011110111100000000000000101",	-- 10581: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 10582: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000010",	-- 10583: 	lli	%r2, 2
"00101000001000100000000000100110",	-- 10584: 	bneq	%r1, %r2, bneq_else.9283
"00111011110000010000000000000011",	-- 10585: 	lw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 10586: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 10587: 	addi	%sp, %sp, 5
"01011000000000000000011001111000",	-- 10588: 	jal	o_diffuse.2646
"10101011110111100000000000000101",	-- 10589: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 10590: 	lw	%ra, [%sp + 4]
"00010100000000010000000000000000",	-- 10591: 	llif	%f1, 1.000000
"00010000000000010011111110000000",	-- 10592: 	lhif	%f1, 1.000000
"00111111111111100000000000000100",	-- 10593: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 10594: 	addi	%sp, %sp, 5
"01011000000000000000010011110001",	-- 10595: 	jal	fless.2532
"10101011110111100000000000000101",	-- 10596: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 10597: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000000",	-- 10598: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 10599: 	bneq	%r1, %r2, bneq_else.9284
"01001111111000000000000000000000",	-- 10600: 	jr	%ra
	-- bneq_else.9284:
"00111011110000010000000000000011",	-- 10601: 	lw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 10602: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 10603: 	addi	%sp, %sp, 5
"01011000000000000000011001010000",	-- 10604: 	jal	o_form.2624
"10101011110111100000000000000101",	-- 10605: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 10606: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000001",	-- 10607: 	lli	%r2, 1
"00101000001000100000000000000110",	-- 10608: 	bneq	%r1, %r2, bneq_else.9286
"00111011110000010000000000000001",	-- 10609: 	lw	%r1, [%sp + 1]
"00111011110000100000000000000011",	-- 10610: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000010",	-- 10611: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 10612: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10613: 	jr	%r26
	-- bneq_else.9286:
"11001100000000100000000000000010",	-- 10614: 	lli	%r2, 2
"00101000001000100000000000000110",	-- 10615: 	bneq	%r1, %r2, bneq_else.9287
"00111011110000010000000000000001",	-- 10616: 	lw	%r1, [%sp + 1]
"00111011110000100000000000000011",	-- 10617: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000000",	-- 10618: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10619: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10620: 	jr	%r26
	-- bneq_else.9287:
"01001111111000000000000000000000",	-- 10621: 	jr	%ra
	-- bneq_else.9283:
"01001111111000000000000000000000",	-- 10622: 	jr	%ra
	-- bgt_else.9282:
"01001111111000000000000000000000",	-- 10623: 	jr	%ra
	-- rt.3049:
"00111011011000110000000000001110",	-- 10624: 	lw	%r3, [%r27 + 14]
"00111011011001000000000000001101",	-- 10625: 	lw	%r4, [%r27 + 13]
"00111011011001010000000000001100",	-- 10626: 	lw	%r5, [%r27 + 12]
"00111011011001100000000000001011",	-- 10627: 	lw	%r6, [%r27 + 11]
"00111011011001110000000000001010",	-- 10628: 	lw	%r7, [%r27 + 10]
"00111011011010000000000000001001",	-- 10629: 	lw	%r8, [%r27 + 9]
"00111011011010010000000000001000",	-- 10630: 	lw	%r9, [%r27 + 8]
"00111011011010100000000000000111",	-- 10631: 	lw	%r10, [%r27 + 7]
"00111011011010110000000000000110",	-- 10632: 	lw	%r11, [%r27 + 6]
"00111011011011000000000000000101",	-- 10633: 	lw	%r12, [%r27 + 5]
"00111011011011010000000000000100",	-- 10634: 	lw	%r13, [%r27 + 4]
"00111011011011100000000000000011",	-- 10635: 	lw	%r14, [%r27 + 3]
"00111011011011110000000000000010",	-- 10636: 	lw	%r15, [%r27 + 2]
"00111011011100000000000000000001",	-- 10637: 	lw	%r16, [%r27 + 1]
"11001100000100010000000000000000",	-- 10638: 	lli	%r17, 0
"10000101110100011000100000000000",	-- 10639: 	add	%r17, %r14, %r17
"00111100001100010000000000000000",	-- 10640: 	sw	%r1, [%r17 + 0]
"11001100000100010000000000000001",	-- 10641: 	lli	%r17, 1
"10000101110100010111000000000000",	-- 10642: 	add	%r14, %r14, %r17
"00111100010011100000000000000000",	-- 10643: 	sw	%r2, [%r14 + 0]
"11001100000011100000000000000000",	-- 10644: 	lli	%r14, 0
"01000000001100010000000000000001",	-- 10645: 	sra	%r17, %r1, 1
"10000101111011100111000000000000",	-- 10646: 	add	%r14, %r15, %r14
"00111110001011100000000000000000",	-- 10647: 	sw	%r17, [%r14 + 0]
"11001100000011100000000000000001",	-- 10648: 	lli	%r14, 1
"01000000010000100000000000000001",	-- 10649: 	sra	%r2, %r2, 1
"10000101111011100111000000000000",	-- 10650: 	add	%r14, %r15, %r14
"00111100010011100000000000000000",	-- 10651: 	sw	%r2, [%r14 + 0]
"11001100000000100000000000000000",	-- 10652: 	lli	%r2, 0
"00010100000000000000000000000000",	-- 10653: 	llif	%f0, 128.000000
"00010000000000000100001100000000",	-- 10654: 	lhif	%f0, 128.000000
"00111100111111100000000000000000",	-- 10655: 	sw	%r7, [%sp + 0]
"00111101001111100000000000000001",	-- 10656: 	sw	%r9, [%sp + 1]
"00111100100111100000000000000010",	-- 10657: 	sw	%r4, [%sp + 2]
"00111101010111100000000000000011",	-- 10658: 	sw	%r10, [%sp + 3]
"00111100101111100000000000000100",	-- 10659: 	sw	%r5, [%sp + 4]
"00111101100111100000000000000101",	-- 10660: 	sw	%r12, [%sp + 5]
"00111101011111100000000000000110",	-- 10661: 	sw	%r11, [%sp + 6]
"00111101101111100000000000000111",	-- 10662: 	sw	%r13, [%sp + 7]
"00111100011111100000000000001000",	-- 10663: 	sw	%r3, [%sp + 8]
"00111101000111100000000000001001",	-- 10664: 	sw	%r8, [%sp + 9]
"00111110000111100000000000001010",	-- 10665: 	sw	%r16, [%sp + 10]
"00111100010111100000000000001011",	-- 10666: 	sw	%r2, [%sp + 11]
"00111100110111100000000000001100",	-- 10667: 	sw	%r6, [%sp + 12]
"10110000000111100000000000001101",	-- 10668: 	sf	%f0, [%sp + 13]
"00111111111111100000000000001110",	-- 10669: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 10670: 	addi	%sp, %sp, 15
"01011000000000000010101000101010",	-- 10671: 	jal	yj_float_of_int
"10101011110111100000000000001111",	-- 10672: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 10673: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001101",	-- 10674: 	lf	%f1, [%sp + 13]
"11101100001000000000000000000000",	-- 10675: 	divf	%f0, %f1, %f0
"00111011110000010000000000001011",	-- 10676: 	lw	%r1, [%sp + 11]
"00111011110000100000000000001100",	-- 10677: 	lw	%r2, [%sp + 12]
"10000100010000010000100000000000",	-- 10678: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 10679: 	sf	%f0, [%r1 + 0]
"00111011110110110000000000001010",	-- 10680: 	lw	%r27, [%sp + 10]
"00111111111111100000000000001110",	-- 10681: 	sw	%ra, [%sp + 14]
"00111011011110100000000000000000",	-- 10682: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001111",	-- 10683: 	addi	%sp, %sp, 15
"01010011010000000000000000000000",	-- 10684: 	jalr	%r26
"10101011110111100000000000001111",	-- 10685: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 10686: 	lw	%ra, [%sp + 14]
"00111011110110110000000000001010",	-- 10687: 	lw	%r27, [%sp + 10]
"00111100001111100000000000001110",	-- 10688: 	sw	%r1, [%sp + 14]
"00111111111111100000000000001111",	-- 10689: 	sw	%ra, [%sp + 15]
"00111011011110100000000000000000",	-- 10690: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010000",	-- 10691: 	addi	%sp, %sp, 16
"01010011010000000000000000000000",	-- 10692: 	jalr	%r26
"10101011110111100000000000010000",	-- 10693: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 10694: 	lw	%ra, [%sp + 15]
"00111011110110110000000000001010",	-- 10695: 	lw	%r27, [%sp + 10]
"00111100001111100000000000001111",	-- 10696: 	sw	%r1, [%sp + 15]
"00111111111111100000000000010000",	-- 10697: 	sw	%ra, [%sp + 16]
"00111011011110100000000000000000",	-- 10698: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010001",	-- 10699: 	addi	%sp, %sp, 17
"01010011010000000000000000000000",	-- 10700: 	jalr	%r26
"10101011110111100000000000010001",	-- 10701: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 10702: 	lw	%ra, [%sp + 16]
"00111011110110110000000000001001",	-- 10703: 	lw	%r27, [%sp + 9]
"00111100001111100000000000010000",	-- 10704: 	sw	%r1, [%sp + 16]
"00111111111111100000000000010001",	-- 10705: 	sw	%ra, [%sp + 17]
"00111011011110100000000000000000",	-- 10706: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010010",	-- 10707: 	addi	%sp, %sp, 18
"01010011010000000000000000000000",	-- 10708: 	jalr	%r26
"10101011110111100000000000010010",	-- 10709: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10710: 	lw	%ra, [%sp + 17]
"00111011110110110000000000001000",	-- 10711: 	lw	%r27, [%sp + 8]
"00111111111111100000000000010001",	-- 10712: 	sw	%ra, [%sp + 17]
"00111011011110100000000000000000",	-- 10713: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010010",	-- 10714: 	addi	%sp, %sp, 18
"01010011010000000000000000000000",	-- 10715: 	jalr	%r26
"10101011110111100000000000010010",	-- 10716: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10717: 	lw	%ra, [%sp + 17]
"00111011110110110000000000000111",	-- 10718: 	lw	%r27, [%sp + 7]
"00111111111111100000000000010001",	-- 10719: 	sw	%ra, [%sp + 17]
"00111011011110100000000000000000",	-- 10720: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010010",	-- 10721: 	addi	%sp, %sp, 18
"01010011010000000000000000000000",	-- 10722: 	jalr	%r26
"10101011110111100000000000010010",	-- 10723: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10724: 	lw	%ra, [%sp + 17]
"00111011110000010000000000000110",	-- 10725: 	lw	%r1, [%sp + 6]
"00111111111111100000000000010001",	-- 10726: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 10727: 	addi	%sp, %sp, 18
"01011000000000000000011010111010",	-- 10728: 	jal	d_vec.2683
"10101011110111100000000000010010",	-- 10729: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10730: 	lw	%ra, [%sp + 17]
"00111011110000100000000000000101",	-- 10731: 	lw	%r2, [%sp + 5]
"00111111111111100000000000010001",	-- 10732: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 10733: 	addi	%sp, %sp, 18
"01011000000000000000010100111011",	-- 10734: 	jal	veccpy.2586
"10101011110111100000000000010010",	-- 10735: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10736: 	lw	%ra, [%sp + 17]
"00111011110000010000000000000110",	-- 10737: 	lw	%r1, [%sp + 6]
"00111011110110110000000000000100",	-- 10738: 	lw	%r27, [%sp + 4]
"00111111111111100000000000010001",	-- 10739: 	sw	%ra, [%sp + 17]
"00111011011110100000000000000000",	-- 10740: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010010",	-- 10741: 	addi	%sp, %sp, 18
"01010011010000000000000000000000",	-- 10742: 	jalr	%r26
"10101011110111100000000000010010",	-- 10743: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10744: 	lw	%ra, [%sp + 17]
"11001100000000010000000000000000",	-- 10745: 	lli	%r1, 0
"00111011110000100000000000000011",	-- 10746: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 10747: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 10748: 	lw	%r1, [%r1 + 0]
"11001100000000100000000000000001",	-- 10749: 	lli	%r2, 1
"10001000001000100000100000000000",	-- 10750: 	sub	%r1, %r1, %r2
"00111011110110110000000000000010",	-- 10751: 	lw	%r27, [%sp + 2]
"00111111111111100000000000010001",	-- 10752: 	sw	%ra, [%sp + 17]
"00111011011110100000000000000000",	-- 10753: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010010",	-- 10754: 	addi	%sp, %sp, 18
"01010011010000000000000000000000",	-- 10755: 	jalr	%r26
"10101011110111100000000000010010",	-- 10756: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10757: 	lw	%ra, [%sp + 17]
"11001100000000100000000000000000",	-- 10758: 	lli	%r2, 0
"11001100000000110000000000000000",	-- 10759: 	lli	%r3, 0
"00111011110000010000000000001111",	-- 10760: 	lw	%r1, [%sp + 15]
"00111011110110110000000000000001",	-- 10761: 	lw	%r27, [%sp + 1]
"00111111111111100000000000010001",	-- 10762: 	sw	%ra, [%sp + 17]
"00111011011110100000000000000000",	-- 10763: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010010",	-- 10764: 	addi	%sp, %sp, 18
"01010011010000000000000000000000",	-- 10765: 	jalr	%r26
"10101011110111100000000000010010",	-- 10766: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10767: 	lw	%ra, [%sp + 17]
"11001100000000010000000000000000",	-- 10768: 	lli	%r1, 0
"11001100000001010000000000000010",	-- 10769: 	lli	%r5, 2
"00111011110000100000000000001110",	-- 10770: 	lw	%r2, [%sp + 14]
"00111011110000110000000000001111",	-- 10771: 	lw	%r3, [%sp + 15]
"00111011110001000000000000010000",	-- 10772: 	lw	%r4, [%sp + 16]
"00111011110110110000000000000000",	-- 10773: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10774: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10775: 	jr	%r26
	-- yj_print_char:
"11010000001000000000000000000000",	-- 10776: 	sendc	%r1
"01001111111000000000000000000000",	-- 10777: 	jr	%ra
	-- yj_create_array:
"11001100000000110000000000000000",	-- 10778: 	lli	%r3, 0
	-- yj_create.loop:
"10000111101000110010000000000000",	-- 10779: 	add	%r4, %hp, %r3
"00111100010001000000000000000000",	-- 10780: 	sw	%r2, [%r4 + 0]
"10100100011000110000000000000001",	-- 10781: 	addi	%r3, %r3, 1
"00110000001000111111111111111101",	-- 10782: 	bgt	%r1, %r3, yj_create.loop
"10000100000111010000100000000000",	-- 10783: 	add	%r1, %r0, %hp
"10000111101000111110100000000000",	-- 10784: 	add	%hp, %hp, %r3
"01001111111000000000000000000000",	-- 10785: 	jr	%ra
	-- yj_create_float_array:
"11001100000000110000000000000000",	-- 10786: 	lli	%r3, 0
	-- yj_create_float.loop:
"10000111101000110010000000000000",	-- 10787: 	add	%r4, %hp, %r3
"10110000000001000000000000000000",	-- 10788: 	sf	%f0, [%r4 + 0]
"10100100011000110000000000000001",	-- 10789: 	addi	%r3, %r3, 1
"00110000001000111111111111111101",	-- 10790: 	bgt	%r1, %r3, yj_create_float.loop
"10000100000111010000100000000000",	-- 10791: 	add	%r1, %r0, %hp
"10000111101000111110100000000000",	-- 10792: 	add	%hp, %hp, %r3
"01001111111000000000000000000000",	-- 10793: 	jr	%ra
	-- yj_float_of_int:
"01100000001000000000000000000000",	-- 10794: 	itof	%f0, %r1
"01001111111000000000000000000000",	-- 10795: 	jr	%ra
	-- yj_int_of_float:
"01100100000000010000000000000000",	-- 10796: 	ftoi	%r1, %f0
"01001111111000000000000000000000",	-- 10797: 	jr	%ra
	-- yj_sqrt:
"11110000000000000000000000000000",	-- 10798: 	sqrt	%f0, %f0
"01001111111000000000000000000000",	-- 10799: 	jr	%ra
	-- yj_floor:
"11110100000000000000000000000000",	-- 10800: 	floor	%f0, %f0
"01001111111000000000000000000000",	-- 10801: 	jr	%ra
	-- yj_read_int:
"11001100000000010000000000000000",	-- 10802: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 10803: 	lli	%r2, 0
"11000100000000010000000000000000",	-- 10804: 	recv	%r1
"01001000001000010000000000001000",	-- 10805: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 10806: 	recv	%r2
"10011100001000100000100000000000",	-- 10807: 	xor	%r1, %r1, %r2
"01001000001000010000000000001000",	-- 10808: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 10809: 	recv	%r2
"10011100001000100000100000000000",	-- 10810: 	xor	%r1, %r1, %r2
"01001000001000010000000000001000",	-- 10811: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 10812: 	recv	%r2
"10011100001000100000100000000000",	-- 10813: 	xor	%r1, %r1, %r2
"01001111111000000000000000000000",	-- 10814: 	jr	%ra
	-- yj_read_float:
"11001100000000010000000000000000",	-- 10815: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 10816: 	lli	%r2, 0
"11000100000000010000000000000000",	-- 10817: 	recv	%r1
"01001000001000010000000000001000",	-- 10818: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 10819: 	recv	%r2
"10011100001000100000100000000000",	-- 10820: 	xor	%r1, %r1, %r2
"01001000001000010000000000001000",	-- 10821: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 10822: 	recv	%r2
"10011100001000100000100000000000",	-- 10823: 	xor	%r1, %r1, %r2
"01001000001000010000000000001000",	-- 10824: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 10825: 	recv	%r2
"10011100001000100000100000000000",	-- 10826: 	xor	%r1, %r1, %r2
"01111100001000000000000000000000",	-- 10827: 	movi2f	%f0, %r1
"01001111111000000000000000000000",	-- 10828: 	jr	%ra
	-- yj_fabs:
"11111000000000000000000000000000",	-- 10829: 	absf	%f0, %f0
"01001111111000000000000000000000",	-- 10830: 	jr	%ra
	-- yj_fneg:
"00011000000000000000000000000000",	-- 10831: 	negf	%f0, %f0
"01001111111000000000000000000000"	-- 10832: 	jr	%ra
);

signal shortened : std_logic_vector(6 downto 0):=(others=>'0');
begin  -- R_rom
  shortened<=addra(6 downto 0);
    douta<=rom(conv_integer(shortened));
end R_rom;
