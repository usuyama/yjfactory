library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;


entity PROM is

  port (
    clka  : in  std_logic;
--    wea   : in  std_logic_vector(0 downto 0);
    addra : in  std_logic_vector(6 downto 0);
--    dina  : in  std_logic_vector(31 downto 0);
    douta : out std_logic_vector(31 downto 0));

end PROM;

architecture R_rom of PROM is

type rom_type is array (0 to 111) of std_logic_vector(31 downto 0);
  constant rom : rom_type:=(
"11001100000111100000000000000000",
"10100100000111110000000000000101",
"11001100000111011100001101010000",
"11001100000000010000000000000001",
"01010100000000000000000000010001",
"11111100000000000000000000000000",
"11001100000000110000000000001010",
"00110000011000010000000000000110",
"11001100000000110000000000001010",
"10001000001000110000100000000000",
"11001100000000110000000000000001",
"10000100010000110001000000000000",
"01010100000000000000000000000110",
"10000100000000100000100000000000",
"01001111111000000000000000000000",
"11001100000000100000000000000000",
"01010100000000000000000000000110",
"11001100000000100000000000000000",
"00110000010000010000000000011010",
"11001100000000100000000000001010",
"00110000010000010000000000010101",
"00111100001111100000000000000000",
"00111111111111100000000000000001",
"10100111110111100000000000000010",
"01011000000000000000000000001111",
"10101011110111100000000000000010",
"00111011110111110000000000000001",
"00111100001111100000000000000001",
"00111111111111100000000000000010",
"10100111110111100000000000000011",
"01011000000000000000000000010001",
"10101011110111100000000000000011",
"00111011110111110000000000000010",
"11001100000000010000000000001010",
"00111011110000100000000000000001",
"10001100010000010000100000000000",
"00111011110000100000000000000000",
"10001000010000010000100000000000",
"11001100000000100000000000110000",
"10000100001000100000100000000000",
"01010100000000000000000000110111",
"11001100000000100000000000110000",
"10000100001000100000100000000000",
"01010100000000000000000000110111",
"11001100000000100000000000101101",
"00111100001111100000000000000000",
"10000100000000100000100000000000",
"00111111111111100000000000000010",
"10100111110111100000000000000011",
"01011000000000000000000000110111",
"10101011110111100000000000000011",
"00111011110111110000000000000010",
"00111011110000010000000000000000",
"10001000000000010000100000000000",
"01010100000000000000000000010001",
"11010000001000000000000000000000",
"01001111111000000000000000000000",
"11001100000000110000000000000000",
"10000111101000110010000000000000",
"00111100010001000000000000000000",
"10100100011000110000000000000001",
"00110000001000111111111111111101",
"10000100000111010000100000000000",
"10000111101000111110100000000000",
"01001111111000000000000000000000",
"11001100000000110000000000000000",
"10000111101000110010000000000000",
"10110000000001000000000000000000",
"10100100011000110000000000000001",
"00110000001000111111111111111101",
"10000100000111010000100000000000",
"10000111101000111110100000000000",
"01001111111000000000000000000000",
"01100000001000000000000000000000",
"01001111111000000000000000000000",
"01100100000000010000000000000000",
"01001111111000000000000000000000",
"11110000000000000000000000000000",
"01001111111000000000000000000000",
"11110100000000000000000000000000",
"01001111111000000000000000000000",
"11001100000000010000000000000000",
"11001100000000100000000000000000",
"11000100000000010000000000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001111111000000000000000000000",
"11001100000000010000000000000000",
"11001100000000100000000000000000",
"11000100000000010000000000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01111100001000000000000000000000",
"01001111111000000000000000000000",
"11111000000000000000000000000000",
"01001111111000000000000000000000",
"00011000000000000000000000000000",
"01001111111000000000000000000000"

	-- entry:                
);                               
signal read_a : std_logic_vector(6 downto 0);
signal shortened : std_logic_vector(6 downto 0):=(others=>'0');
begin  -- R_rom
  process(clka)
    begin
    if (clka'event and clka='1') then
      read_a<=addra;
    end if;
  end process;
  shortened<=read_a(6 downto 0);
    douta<=rom(conv_integer(shortened));
end R_rom;

















