library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;


entity PROM is

  port (
    clka  : in  std_logic;
--    wea   : in  std_logic_vector(0 downto 0);
    addra : in  std_logic_vector(6 downto 0);
--    dina  : in  std_logic_vector(31 downto 0);
    douta : out std_logic_vector(31 downto 0));

end PROM;

architecture R_rom of PROM is

type rom_type is array (0 to 179) of std_logic_vector(31 downto 0);
  constant rom : rom_type:=(
	-- entry:
"11001100000111100000000000000000",	-- 0: 	lli	%sp, 0
"10100100000111110000000000100010",	-- 1: 	addi	%ra, %r0, halt
"11001100000111011100001101010000",	-- 2: 	lli	%hp, 50000
"00010100000000001100110011001101",	-- 3: 	llif	%f0, 0.100000
"00010000000000000011110111001100",	-- 4: 	lhif	%f0, 0.100000
"00111111111111100000000000000000",	-- 5: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 6: 	addi	%sp, %sp, 1
"01011000000000000000000001011011",	-- 7: 	jal	f.104
"10101011110111100000000000000001",	-- 8: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 9: 	lw	%ra, [%sp + 0]
"00010100000000000000000000000000",	-- 10: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 11: 	lhif	%f0, 1.000000
"00111111111111100000000000000000",	-- 12: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 13: 	addi	%sp, %sp, 1
"01011000000000000000000001011011",	-- 14: 	jal	f.104
"10101011110111100000000000000001",	-- 15: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 16: 	lw	%ra, [%sp + 0]
"00010100000000000000000000000000",	-- 17: 	llif	%f0, 2.000000
"00010000000000000100000000000000",	-- 18: 	lhif	%f0, 2.000000
"00111111111111100000000000000000",	-- 19: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 20: 	addi	%sp, %sp, 1
"01011000000000000000000001011011",	-- 21: 	jal	f.104
"10101011110111100000000000000001",	-- 22: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 23: 	lw	%ra, [%sp + 0]
"00010100000000000000000000000000",	-- 24: 	llif	%f0, 5.000000
"00010000000000000100000010100000",	-- 25: 	lhif	%f0, 5.000000
"00111111111111100000000000000000",	-- 26: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 27: 	addi	%sp, %sp, 1
"01011000000000000000000001011011",	-- 28: 	jal	f.104
"10101011110111100000000000000001",	-- 29: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 30: 	lw	%ra, [%sp + 0]
"00010100000000000000000000000000",	-- 31: 	llif	%f0, 10.000000
"00010000000000000100000100100000",	-- 32: 	lhif	%f0, 10.000000
"01010100000000000000000001011011",	-- 33: 	j	f.104
	-- halt:
"11111100000000000000000000000000",	-- 34: 	halt
	-- atan.102:
"10110000000111100000000000000000",	-- 35: 	sf	%f0, [%sp + 0]
"00111111111111100000000000000001",	-- 36: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 37: 	addi	%sp, %sp, 2
"01011000000000000000000010100101",	-- 38: 	jal	yj_fabs
"10101011110111100000000000000010",	-- 39: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 40: 	lw	%ra, [%sp + 1]
"00010100000000011001100110011010",	-- 41: 	llif	%f1, 0.150000
"00010000000000010011111000011001",	-- 42: 	lhif	%f1, 0.150000
"00100000000000010000000000010011",	-- 43: 	bgtf	%f0, %f1, bgtf_else.246
"10010011110000000000000000000000",	-- 44: 	lf	%f0, [%sp + 0]
"11101000000000000000100000000000",	-- 45: 	mulf	%f1, %f0, %f0
"00010100000000100000000000000000",	-- 46: 	llif	%f2, 1.000000
"00010000000000100011111110000000",	-- 47: 	lhif	%f2, 1.000000
"00010100000000111010101010011111",	-- 48: 	llif	%f3, -0.333333
"00010000000000111011111010101010",	-- 49: 	lhif	%f3, -0.333333
"00010100000001001100110011001101",	-- 50: 	llif	%f4, 0.200000
"00010000000001000011111001001100",	-- 51: 	lhif	%f4, 0.200000
"00010100000001010100100100011011",	-- 52: 	llif	%f5, 0.142857
"00010000000001010011111000010010",	-- 53: 	lhif	%f5, 0.142857
"11101000001001010010100000000000",	-- 54: 	mulf	%f5, %f1, %f5
"11100000100001010010000000000000",	-- 55: 	addf	%f4, %f4, %f5
"11101000001001000010000000000000",	-- 56: 	mulf	%f4, %f1, %f4
"11100000011001000001100000000000",	-- 57: 	addf	%f3, %f3, %f4
"11101000001000110000100000000000",	-- 58: 	mulf	%f1, %f1, %f3
"11100000010000010000100000000000",	-- 59: 	addf	%f1, %f2, %f1
"11101000000000010000000000000000",	-- 60: 	mulf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 61: 	jr	%ra
	-- bgtf_else.246:
"00010100000000000000000000000000",	-- 62: 	llif	%f0, -1.000000
"00010000000000001011111110000000",	-- 63: 	lhif	%f0, -1.000000
"00010100000000010000000000000000",	-- 64: 	llif	%f1, 1.000000
"00010000000000010011111110000000",	-- 65: 	lhif	%f1, 1.000000
"10010011110000100000000000000000",	-- 66: 	lf	%f2, [%sp + 0]
"11101000010000100001100000000000",	-- 67: 	mulf	%f3, %f2, %f2
"11100000001000110000100000000000",	-- 68: 	addf	%f1, %f1, %f3
"10110000000111100000000000000001",	-- 69: 	sf	%f0, [%sp + 1]
"00001100001000000000000000000000",	-- 70: 	movf	%f0, %f1
"00111111111111100000000000000010",	-- 71: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 72: 	addi	%sp, %sp, 3
"01011000000000000000000010000110",	-- 73: 	jal	yj_sqrt
"10101011110111100000000000000011",	-- 74: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 75: 	lw	%ra, [%sp + 2]
"10010011110000010000000000000001",	-- 76: 	lf	%f1, [%sp + 1]
"11100000001000000000000000000000",	-- 77: 	addf	%f0, %f1, %f0
"10010011110000010000000000000000",	-- 78: 	lf	%f1, [%sp + 0]
"11101100000000010000000000000000",	-- 79: 	divf	%f0, %f0, %f1
"00010100000000010000000000000000",	-- 80: 	llif	%f1, 2.000000
"00010000000000010100000000000000",	-- 81: 	lhif	%f1, 2.000000
"10110000001111100000000000000010",	-- 82: 	sf	%f1, [%sp + 2]
"00111111111111100000000000000011",	-- 83: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 84: 	addi	%sp, %sp, 4
"01011000000000000000000000100011",	-- 85: 	jal	atan.102
"10101011110111100000000000000100",	-- 86: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 87: 	lw	%ra, [%sp + 3]
"10010011110000010000000000000010",	-- 88: 	lf	%f1, [%sp + 2]
"11101000001000000000000000000000",	-- 89: 	mulf	%f0, %f1, %f0
"01001111111000000000000000000000",	-- 90: 	jr	%ra
	-- f.104:
"10110000000111100000000000000000",	-- 91: 	sf	%f0, [%sp + 0]
"00111111111111100000000000000001",	-- 92: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 93: 	addi	%sp, %sp, 2
"01011000000000000000000000100011",	-- 94: 	jal	atan.102
"10101011110111100000000000000010",	-- 95: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 96: 	lw	%ra, [%sp + 1]
"00111111111111100000000000000001",	-- 97: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 98: 	addi	%sp, %sp, 2
"01011000000000000000000010101001",	-- 99: 	jal	yj_print_float_binary
"10101011110111100000000000000010",	-- 100: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 101: 	lw	%ra, [%sp + 1]
"00010100000000000000000000000000",	-- 102: 	llif	%f0, -1.000000
"00010000000000001011111110000000",	-- 103: 	lhif	%f0, -1.000000
"10010011110000010000000000000000",	-- 104: 	lf	%f1, [%sp + 0]
"11101000000000010000000000000000",	-- 105: 	mulf	%f0, %f0, %f1
"00111111111111100000000000000001",	-- 106: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 107: 	addi	%sp, %sp, 2
"01011000000000000000000000100011",	-- 108: 	jal	atan.102
"10101011110111100000000000000010",	-- 109: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 110: 	lw	%ra, [%sp + 1]
"01010100000000000000000010101001",	-- 111: 	j	yj_print_float_binary
	-- yj_print_char:
"11010000001000000000000000000000",	-- 112: 	sendc	%r1
"01001111111000000000000000000000",	-- 113: 	jr	%ra
	-- yj_create_array:
"11001100000000110000000000000000",	-- 114: 	lli	%r3, 0
	-- yj_create.loop:
"10000111101000110010000000000000",	-- 115: 	add	%r4, %hp, %r3
"00111100010001000000000000000000",	-- 116: 	sw	%r2, [%r4 + 0]
"10100100011000110000000000000001",	-- 117: 	addi	%r3, %r3, 1
"00110000001000111111111111111101",	-- 118: 	bgt	%r1, %r3, yj_create.loop
"10000100000111010000100000000000",	-- 119: 	add	%r1, %r0, %hp
"10000111101000111110100000000000",	-- 120: 	add	%hp, %hp, %r3
"01001111111000000000000000000000",	-- 121: 	jr	%ra
	-- yj_create_float_array:
"11001100000000110000000000000000",	-- 122: 	lli	%r3, 0
	-- yj_create_float.loop:
"10000111101000110010000000000000",	-- 123: 	add	%r4, %hp, %r3
"10110000000001000000000000000000",	-- 124: 	sf	%f0, [%r4 + 0]
"10100100011000110000000000000001",	-- 125: 	addi	%r3, %r3, 1
"00110000001000111111111111111101",	-- 126: 	bgt	%r1, %r3, yj_create_float.loop
"10000100000111010000100000000000",	-- 127: 	add	%r1, %r0, %hp
"10000111101000111110100000000000",	-- 128: 	add	%hp, %hp, %r3
"01001111111000000000000000000000",	-- 129: 	jr	%ra
	-- yj_float_of_int:
"01100000001000000000000000000000",	-- 130: 	itof	%f0, %r1
"01001111111000000000000000000000",	-- 131: 	jr	%ra
	-- yj_int_of_float:
"01100100000000010000000000000000",	-- 132: 	ftoi	%r1, %f0
"01001111111000000000000000000000",	-- 133: 	jr	%ra
	-- yj_sqrt:
"11110000000000000000000000000000",	-- 134: 	sqrt	%f0, %f0
"01001111111000000000000000000000",	-- 135: 	jr	%ra
	-- yj_floor:
"11110100000000000000000000000000",	-- 136: 	floor	%f0, %f0
"01001111111000000000000000000000",	-- 137: 	jr	%ra
	-- yj_read_int:
"11001100000000010000000000000000",	-- 138: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 139: 	lli	%r2, 0
"11000100000000010000000000000000",	-- 140: 	recv	%r1
"01001000001000010000000000001000",	-- 141: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 142: 	recv	%r2
"10011100001000100000100000000000",	-- 143: 	xor	%r1, %r1, %r2
"01001000001000010000000000001000",	-- 144: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 145: 	recv	%r2
"10011100001000100000100000000000",	-- 146: 	xor	%r1, %r1, %r2
"01001000001000010000000000001000",	-- 147: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 148: 	recv	%r2
"10011100001000100000100000000000",	-- 149: 	xor	%r1, %r1, %r2
"01001111111000000000000000000000",	-- 150: 	jr	%ra
	-- yj_read_float:
"11001100000000010000000000000000",	-- 151: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 152: 	lli	%r2, 0
"11000100000000010000000000000000",	-- 153: 	recv	%r1
"01001000001000010000000000001000",	-- 154: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 155: 	recv	%r2
"10011100001000100000100000000000",	-- 156: 	xor	%r1, %r1, %r2
"01001000001000010000000000001000",	-- 157: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 158: 	recv	%r2
"10011100001000100000100000000000",	-- 159: 	xor	%r1, %r1, %r2
"01001000001000010000000000001000",	-- 160: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 161: 	recv	%r2
"10011100001000100000100000000000",	-- 162: 	xor	%r1, %r1, %r2
"01111100001000000000000000000000",	-- 163: 	movi2f	%f0, %r1
"01001111111000000000000000000000",	-- 164: 	jr	%ra
	-- yj_fabs:
"11111000000000000000000000000000",	-- 165: 	absf	%f0, %f0
"01001111111000000000000000000000",	-- 166: 	jr	%ra
	-- yj_fneg:
"00011000000000000000000000000000",	-- 167: 	negf	%f0, %f0
"01001111111000000000000000000000",	-- 168: 	jr	%ra
	-- yj_print_float_binary:
"01011100000000010000000000000000",	-- 169: 	movf2i	%r1, %f0
"11010000001000000000000000000000",	-- 170: 	sendc	%r1
"01000000001000010000000000001000",	-- 171: 	sra	%r1, %r1, 8
"11010000001000000000000000000000",	-- 172: 	sendc	%r1
"01000000001000010000000000001000",	-- 173: 	sra	%r1, %r1, 8
"11010000001000000000000000000000",	-- 174: 	sendc	%r1
"01000000001000010000000000001000",	-- 175: 	sra	%r1, %r1, 8
"11010000001000000000000000000000",	-- 176: 	sendc	%r1
"11001100000000010000000000001010",	-- 177: 	lli	%r1, 10
"11010000001000000000000000000000",	-- 178: 	sendc	%r1
"01001111111000000000000000000000"	-- 179: 	jr	%ra
);

signal shortened : std_logic_vector(6 downto 0):=(others=>'0');
begin  -- R_rom
  shortened<=addra(6 downto 0);
    douta<=rom(conv_integer(shortened));
end R_rom;
