library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;


entity PROM is
  
  port (
    clka  : in  std_logic;
--    wea   : in  std_logic_vector(0 downto 0);
    addra : in  std_logic_vector(31 downto 0);
--    dina  : in  std_logic_vector(31 downto 0);
    douta : out std_logic_vector(31 downto 0));

end PROM;

architecture R_rom of PROM is
type rom_type is array (0 to 34) of std_logic_vector(31 downto 0);
constant rom : rom_type:=(
"11001000000111100000000000000000",     --0
"11001000000111110000000000000000",     --1
"11001000000111010010011100010000",     --2
"11001000000000010000000000000101",     --3
"00111111111111100000000000000000",     --4
"10100111110111100000000000000001",     --5
"01011000000000000000000000001010",     --6
"10101011110111100000000000000001",     --7
"00111011110111110000000000000000",     --8
"11000000000000000000000000000000",     --9
"11001000000000100000000000000001",     --10
"00110000001000100000000000000010",     --11
"01001111111000000000000000000000",     --12
"11001000000000100000000000000001",     --13
"10001000001000100001000000000000",     --14
"00111100001111100000000000000000",     --15
"10000100000000100000100000000000",     --10
"00111111111111100000000000000001",     --11
"10100111110111100000000000000010",     --12
"01011000000000000000000000001010",     --13
"10101011110111100000000000000010",     --14
"00111011110111110000000000000001",     --15
"11001000000000100000000000000010",     --16
"00111011110000110000000000000000",     --17
"10001000011000100001000000000000",     --18
"00111100001111100000000000000001",     --19
"10000100000000100000100000000000",     --1a
"00111111111111100000000000000010",     --1b
"10100111110111100000000000000011",     --1c
"01011000000000000000000000001010",     --1d
"10101011110111100000000000000011",     --1e
"00111011110111110000000000000010",     --1f
"00111011110000100000000000000001",     --20
"10000100010000010000100000000000",     --21
"01001111111000000000000000000000"      --22
--"00000000000000000000000000000000",
--"10100100001000010000000000001010",
--"00111100001000010000000000000000",
--"00111000001000100000000000000000",
--"10000100010000010001100000000000" 

);

signal shortened : std_logic_vector(5 downto 0):=(others=>'0');
  
begin  -- R_rom
  shortened<=addra(5 downto 0);
    douta<=rom(conv_integer(shortened));
end R_rom;







