library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;


entity PROM is

  port (
    clka  : in  std_logic;
--    wea   : in  std_logic_vector(0 downto 0);
    addra : in  std_logic_vector(6 downto 0);
--    dina  : in  std_logic_vector(31 downto 0);
    douta : out std_logic_vector(31 downto 0));

end PROM;

architecture R_rom of PROM is
-- %r1 = 9169 expected
type rom_type is array (0 to 78) of std_logic_vector(31 downto 0);
  constant rom : rom_type:=(
	-- entry:
"11001100000111100000000000000000",	-- 1: 	lli	%sp, 0
"10100100000111110000000000001000",	-- 2: 	addi	%ra, %r0, halt
"11001100000111011100001101010000",	-- 3: 	lli	%hp, 50000
"11001100000000010000000000000011",	-- 4: 	lli	%r1, 3
"11001100000000100000000000000011",	-- 5: 	lli	%r2, 3
"11001100000000110000000000000000",	-- 6: 	lli	%r3, 0
"11001100000001000000000000000000",	-- 7: 	lli	%r4, 0
"01010100000000000000000000001001",	-- 8: 	j	f.130
	-- halt:
"11111100000000000000000000000000",	-- 9: 	halt
	-- f.130:
"11001100000001010000000001100100",	-- 10: 	lli	%r5, 100
"00110000011001010000000000100111",	-- 11: 	bgt	%r3, %r5, bgt_else.295
"11001100000001010010011100010000",	-- 12: 	lli	%r5, 10000
"00110000010001010000000000011110",	-- 13: 	bgt	%r2, %r5, bgt_else.296
"11001100000001010010011100010000",	-- 14: 	lli	%r5, 10000
"00110000001001010000000000010010",	-- 15: 	bgt	%r1, %r5, bgt_else.297
"00110000010000010000000000001001",	-- 16: 	bgt	%r2, %r1, bgt_else.298
"10001100001000100010100000000000",	-- 17: 	mul	%r5, %r1, %r2
"10000100010000010001000000000000",	-- 18: 	add	%r2, %r2, %r1
"11001100000000010000000000000001",	-- 19: 	lli	%r1, 1
"10000100011000010001100000000000",	-- 20: 	add	%r3, %r3, %r1
"11001100000000010000000000000001",	-- 21: 	lli	%r1, 1
"10001000100000010010000000000000",	-- 22: 	sub	%r4, %r4, %r1
"10000100000001010000100000000000",	-- 23: 	add	%r1, %r0, %r5
"01010100000000000000000000001001",	-- 24: 	j	f.130
	-- bgt_else.298:
"10001100001000100010100000000000",	-- 25: 	mul	%r5, %r1, %r2
"10001000010000010001000000000000",	-- 26: 	sub	%r2, %r2, %r1
"11001100000000010000000000000001",	-- 27: 	lli	%r1, 1
"10000100011000010001100000000000",	-- 28: 	add	%r3, %r3, %r1
"11001100000000010000000000000001",	-- 29: 	lli	%r1, 1
"10001000100000010010000000000000",	-- 30: 	sub	%r4, %r4, %r1
"10000100000001010000100000000000",	-- 31: 	add	%r1, %r0, %r5
"01010100000000000000000000001001",	-- 32: 	j	f.130
	-- bgt_else.297:
"10001100001000100001000000000000",	-- 33: 	mul	%r2, %r1, %r2
"01000000001000010000000000000001",	-- 34: 	sra	%r1, %r1, 1
"11001100000001010000000000000001",	-- 35: 	lli	%r5, 1
"10000100011001010001100000000000",	-- 36: 	add	%r3, %r3, %r5
"11001100000001010000000000000001",	-- 37: 	lli	%r5, 1
"10001000100001010010000000000000",	-- 38: 	sub	%r4, %r4, %r5
"10000100000000101101000000000000",	-- 39: 	add	%r26, %r0, %r2
"10000100000000010001000000000000",	-- 40: 	add	%r2, %r0, %r1
"10000100000110100000100000000000",	-- 41: 	add	%r1, %r0, %r26
"01010100000000000000000000001001",	-- 42: 	j	f.130
	-- bgt_else.296:
"10001100001000100000100000000000",	-- 43: 	mul	%r1, %r1, %r2
"01000000010000100000000000000001",	-- 44: 	sra	%r2, %r2, 1
"11001100000001010000000000000001",	-- 45: 	lli	%r5, 1
"10000100011001010001100000000000",	-- 46: 	add	%r3, %r3, %r5
"11001100000001010000000000000001",	-- 47: 	lli	%r5, 1
"10001000100001010010000000000000",	-- 48: 	sub	%r4, %r4, %r5
"01010100000000000000000000001001",	-- 49: 	j	f.130
	-- bgt_else.295:
"11001100000001010000000001100101",	-- 50: 	lli	%r5, 101
"00110000011001010000000000011010",	-- 51: 	bgt	%r3, %r5, bgt_else.299
"11001100000001011111111110011100",	-- 52: 	lli	%r5, -100
"11001000000001011111111111111111",	-- 53: 	lhi	%r5, -100
"00110000101001000000000000000100",	-- 54: 	bgt	%r5, %r4, bgt_else.300
"11001100000000011111111111111100",	-- 55: 	lli	%r1, -4
"11001000000000011111111111111111",	-- 56: 	lhi	%r1, -4
"01001111111000000000000000000000",	-- 57: 	jr	%ra
	-- bgt_else.300:
"11001100000001011111111110011011",	-- 58: 	lli	%r5, -101
"11001000000001011111111111111111",	-- 59: 	lhi	%r5, -101
"00110000101001000000000000001110",	-- 60: 	bgt	%r5, %r4, bgt_else.301
"11001100000001010000000001100101",	-- 61: 	lli	%r5, 101
"00101000011001010000000000001001",	-- 62: 	bneq	%r3, %r5, bneq_else.302
"11001100000000111111111110011011",	-- 63: 	lli	%r3, -101
"11001000000000111111111111111111",	-- 64: 	lhi	%r3, -101
"00101000100000110000000000000011",	-- 65: 	bneq	%r4, %r3, bneq_else.303
"10000100001000100000100000000000",	-- 66: 	add	%r1, %r1, %r2
"01001111111000000000000000000000",	-- 67: 	jr	%ra
	-- bneq_else.303:
"11001100000000011111111111111111",	-- 68: 	lli	%r1, -1
"11001000000000011111111111111111",	-- 69: 	lhi	%r1, -1
"01001111111000000000000000000000",	-- 70: 	jr	%ra
	-- bneq_else.302:
"11001100000000011111111111111110",	-- 71: 	lli	%r1, -2
"11001000000000011111111111111111",	-- 72: 	lhi	%r1, -2
"01001111111000000000000000000000",	-- 73: 	jr	%ra
	-- bgt_else.301:
"11001100000000011111111111111101",	-- 74: 	lli	%r1, -3
"11001000000000011111111111111111",	-- 75: 	lhi	%r1, -3
"01001111111000000000000000000000",	-- 76: 	jr	%ra
	-- bgt_else.299:
"11001100000000011111111111111011",	-- 77: 	lli	%r1, -5
"11001000000000011111111111111111",	-- 78: 	lhi	%r1, -5
"01001111111000000000000000000000"	-- 79: 	jr	%ra
);

signal shortened : std_logic_vector(6 downto 0):=(others=>'0');
begin  -- R_rom
  shortened<=addra(6 downto 0);
    douta<=rom(conv_integer(shortened));
end R_rom;
