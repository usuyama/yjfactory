library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity instmem is
      port(
        CLK : in std_logic;
        BUBBLE: in std_logic;
        ADRS : in std_logic_vector (13 downto 0);
        DOUT:out std_logic_vector(31 downto 0)
    );
end instmem;

architecture behav of instmem is
type RamType is array(0 to 16383) of std_logic_vector(31 downto 0);
signal RAM:RamType :=(
"11001100000111100000000000000000",
"10100100000111110000000000001100",
"11001100000111011100001101010000",
"11001100000000010000000000011110",
"00111111111111100000000000000000",
"10100111110111100000000000000001",
"01011000000000000000000001000011",
"10101011110111100000000000000001",
"00111011110111110000000000000000",
"11001100000000101011001000101000",
"11001000000000100000000000001100",
"01010100000000000000000000111110",
"11111100000000000000000000000000",
"11001100000000110000000000001010",
"00110000011000010000000000000110",
"11001100000000110000000000001010",
"10001000001000110000100000000000",
"11001100000000110000000000000001",
"10000100010000110001000000000000",
"01010100000000000000000000001101",
"10000100000000100000100000000000",
"01001111111000000000000000000000",
"11001100000000100000000000000000",
"01010100000000000000000000001101",
"11001100000000100000000000000000",
"00110000010000010000000000011010",
"11001100000000100000000000001010",
"00110000010000010000000000010101",
"00111100001111100000000000000000",
"00111111111111100000000000000001",
"10100111110111100000000000000010",
"01011000000000000000000000010110",
"10101011110111100000000000000010",
"00111011110111110000000000000001",
"00111100001111100000000000000001",
"00111111111111100000000000000010",
"10100111110111100000000000000011",
"01011000000000000000000000011000",
"10101011110111100000000000000011",
"00111011110111110000000000000010",
"11001100000000010000000000001010",
"00111011110000100000000000000001",
"10001100010000010000100000000000",
"00111011110000100000000000000000",
"10001000010000010000100000000000",
"11001100000000100000000000110000",
"10000100001000100000100000000000",
"01010100000000000000000001011100",
"11001100000000100000000000110000",
"10000100001000100000100000000000",
"01010100000000000000000001011100",
"11001100000000100000000000101101",
"00111100001111100000000000000000",
"10000100000000100000100000000000",
"00111111111111100000000000000010",
"10100111110111100000000000000011",
"01011000000000000000000001011100",
"10101011110111100000000000000011",
"00111011110111110000000000000010",
"00111011110000010000000000000000",
"10001000000000010000100000000000",
"01010100000000000000000000011000",
"00101000001000100000000000000011",
"11001100000000010000000000000001",
"01010100000000000000000000011000",
"11001100000000010000000000000000",
"01010100000000000000000000011000",
"11001100000000100000000000000001",
"00110000001000100000000000000010",
"01001111111000000000000000000000",
"11001100000000100000000000000001",
"10001000001000100001000000000000",
"00111100001111100000000000000000",
"10000100000000100000100000000000",
"00111111111111100000000000000001",
"10100111110111100000000000000010",
"01011000000000000000000001000011",
"10101011110111100000000000000010",
"00111011110111110000000000000001",
"11001100000000100000000000000010",
"00111011110000110000000000000000",
"10001000011000100001000000000000",
"00111100001111100000000000000001",
"10000100000000100000100000000000",
"00111111111111100000000000000010",
"10100111110111100000000000000011",
"01011000000000000000000001000011",
"10101011110111100000000000000011",
"00111011110111110000000000000010",
"00111011110000100000000000000001",
"10000100010000010000100000000000",
"01001111111000000000000000000000",
"11010000001000000000000000000000",
"01001111111000000000000000000000",
"11001100000000110000000000000000",
"10000111101000110010000000000000",
"00111100010001000000000000000000",
"10100100011000110000000000000001",
"00110000001000111111111111111101",
"10000100000111010000100000000000",
"10000111101000111110100000000000",
"01001111111000000000000000000000",
"11001100000000110000000000000000",
"10000111101000110010000000000000",
"10110000000001000000000000000000",
"10100100011000110000000000000001",
"00110000001000111111111111111101",
"10000100000111010000100000000000",
"10000111101000111110100000000000",
"01001111111000000000000000000000",
"01100000001000000000000000000000",
"01001111111000000000000000000000",
"01100100000000010000000000000000",
"01001111111000000000000000000000",
"11110000000000000000000000000000",
"01001111111000000000000000000000",
"11110100000000000000000000000000",
"01001111111000000000000000000000",
"11001100000000010000000000000000",
"11001100000000100000000000000000",
"11000100000000010000000000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001111111000000000000000000000",
"11001100000000010000000000000000",
"11001100000000100000000000000000",
"11000100000000010000000000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01001000001000010000000000001000",
"11000100000000100000000000000000",
"10011100001000100000100000000000",
"01111100001000000000000000000000",
"01001111111000000000000000000000",
"11111000000000000000000000000000",
"01001111111000000000000000000000",
"00011000000000000000000000000000",
"01001111111000000000000000000000",
others => (others => '0'));

begin
  process(clk) begin
   if rising_edge(clk) then
     if BUBBLE='1' then
       DOUT <= x"00000000";
     else
       DOUT <= RAM(conv_integer (ADRS));
     end if;
   end if;
  end process;
end behav;
