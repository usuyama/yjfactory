library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;


entity PROM is

  port (
    clka  : in  std_logic;
--    wea   : in  std_logic_vector(0 downto 0);
    addra : in  std_logic_vector(6 downto 0);
--    dina  : in  std_logic_vector(31 downto 0);
    douta : out std_logic_vector(31 downto 0));

end PROM;

architecture R_rom of PROM is

type rom_type is array (0 to 10834) of std_logic_vector(31 downto 0);
  constant rom : rom_type:=(
	-- entry:
"00000000000000000000000000000000",	-- 0: 	nop
"11001100000000010000000010101010",	-- 1: 	lli	%r1, 170
"11010000001000000000000000000000",	-- 2: 	sendc	%r1
"11001100000111100000000000000000",	-- 3: 	lli	%sp, 0
"10100100000111110000001111110110",	-- 4: 	addi	%ra, %r0, halt
"11001100000111011100001101010000",	-- 5: 	lli	%hp, 50000
"11001100000000010000000000000001",	-- 6: 	lli	%r1, 1
"11001100000000100000000000000000",	-- 7: 	lli	%r2, 0
"00111111111111100000000000000000",	-- 8: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 9: 	addi	%sp, %sp, 1
"01011000000000000010101000011100",	-- 10: 	jal	yj_create_array
"10101011110111100000000000000001",	-- 11: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 12: 	lw	%ra, [%sp + 0]
"11001100000000100000000000000000",	-- 13: 	lli	%r2, 0
"00010100000000000000000000000000",	-- 14: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 15: 	lhif	%f0, 0.000000
"00111100001111100000000000000000",	-- 16: 	sw	%r1, [%sp + 0]
"10000100000000100000100000000000",	-- 17: 	add	%r1, %r0, %r2
"00111111111111100000000000000001",	-- 18: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 19: 	addi	%sp, %sp, 2
"01011000000000000010101000100100",	-- 20: 	jal	yj_create_float_array
"10101011110111100000000000000010",	-- 21: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 22: 	lw	%ra, [%sp + 1]
"11001100000000100000000000111100",	-- 23: 	lli	%r2, 60
"11001100000000110000000000000000",	-- 24: 	lli	%r3, 0
"11001100000001000000000000000000",	-- 25: 	lli	%r4, 0
"11001100000001010000000000000000",	-- 26: 	lli	%r5, 0
"11001100000001100000000000000000",	-- 27: 	lli	%r6, 0
"11001100000001110000000000000000",	-- 28: 	lli	%r7, 0
"10000100000111010100000000000000",	-- 29: 	add	%r8, %r0, %hp
"10100111101111010000000000001011",	-- 30: 	addi	%hp, %hp, 11
"00111100001010000000000000001010",	-- 31: 	sw	%r1, [%r8 + 10]
"00111100001010000000000000001001",	-- 32: 	sw	%r1, [%r8 + 9]
"00111100001010000000000000001000",	-- 33: 	sw	%r1, [%r8 + 8]
"00111100001010000000000000000111",	-- 34: 	sw	%r1, [%r8 + 7]
"00111100111010000000000000000110",	-- 35: 	sw	%r7, [%r8 + 6]
"00111100001010000000000000000101",	-- 36: 	sw	%r1, [%r8 + 5]
"00111100001010000000000000000100",	-- 37: 	sw	%r1, [%r8 + 4]
"00111100110010000000000000000011",	-- 38: 	sw	%r6, [%r8 + 3]
"00111100101010000000000000000010",	-- 39: 	sw	%r5, [%r8 + 2]
"00111100100010000000000000000001",	-- 40: 	sw	%r4, [%r8 + 1]
"00111100011010000000000000000000",	-- 41: 	sw	%r3, [%r8 + 0]
"10000100000010000000100000000000",	-- 42: 	add	%r1, %r0, %r8
"10000100000000101101000000000000",	-- 43: 	add	%r26, %r0, %r2
"10000100000000010001000000000000",	-- 44: 	add	%r2, %r0, %r1
"10000100000110100000100000000000",	-- 45: 	add	%r1, %r0, %r26
"00111111111111100000000000000001",	-- 46: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 47: 	addi	%sp, %sp, 2
"01011000000000000010101000011100",	-- 48: 	jal	yj_create_array
"10101011110111100000000000000010",	-- 49: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 50: 	lw	%ra, [%sp + 1]
"11001100000000100000000000000011",	-- 51: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 52: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 53: 	lhif	%f0, 0.000000
"00111100001111100000000000000001",	-- 54: 	sw	%r1, [%sp + 1]
"10000100000000100000100000000000",	-- 55: 	add	%r1, %r0, %r2
"00111111111111100000000000000010",	-- 56: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 57: 	addi	%sp, %sp, 3
"01011000000000000010101000100100",	-- 58: 	jal	yj_create_float_array
"10101011110111100000000000000011",	-- 59: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 60: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000011",	-- 61: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 62: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 63: 	lhif	%f0, 0.000000
"00111100001111100000000000000010",	-- 64: 	sw	%r1, [%sp + 2]
"10000100000000100000100000000000",	-- 65: 	add	%r1, %r0, %r2
"00111111111111100000000000000011",	-- 66: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 67: 	addi	%sp, %sp, 4
"01011000000000000010101000100100",	-- 68: 	jal	yj_create_float_array
"10101011110111100000000000000100",	-- 69: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 70: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000011",	-- 71: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 72: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 73: 	lhif	%f0, 0.000000
"00111100001111100000000000000011",	-- 74: 	sw	%r1, [%sp + 3]
"10000100000000100000100000000000",	-- 75: 	add	%r1, %r0, %r2
"00111111111111100000000000000100",	-- 76: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 77: 	addi	%sp, %sp, 5
"01011000000000000010101000100100",	-- 78: 	jal	yj_create_float_array
"10101011110111100000000000000101",	-- 79: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 80: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000001",	-- 81: 	lli	%r2, 1
"00010100000000000000000000000000",	-- 82: 	llif	%f0, 255.000000
"00010000000000000100001101111111",	-- 83: 	lhif	%f0, 255.000000
"00111100001111100000000000000100",	-- 84: 	sw	%r1, [%sp + 4]
"10000100000000100000100000000000",	-- 85: 	add	%r1, %r0, %r2
"00111111111111100000000000000101",	-- 86: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 87: 	addi	%sp, %sp, 6
"01011000000000000010101000100100",	-- 88: 	jal	yj_create_float_array
"10101011110111100000000000000110",	-- 89: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 90: 	lw	%ra, [%sp + 5]
"11001100000000100000000000110010",	-- 91: 	lli	%r2, 50
"11001100000000110000000000000001",	-- 92: 	lli	%r3, 1
"11001100000001001111111111111111",	-- 93: 	lli	%r4, -1
"11001000000001001111111111111111",	-- 94: 	lhi	%r4, -1
"00111100001111100000000000000101",	-- 95: 	sw	%r1, [%sp + 5]
"00111100010111100000000000000110",	-- 96: 	sw	%r2, [%sp + 6]
"10000100000001000001000000000000",	-- 97: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 98: 	add	%r1, %r0, %r3
"00111111111111100000000000000111",	-- 99: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 100: 	addi	%sp, %sp, 8
"01011000000000000010101000011100",	-- 101: 	jal	yj_create_array
"10101011110111100000000000001000",	-- 102: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 103: 	lw	%ra, [%sp + 7]
"10000100000000010001000000000000",	-- 104: 	add	%r2, %r0, %r1
"00111011110000010000000000000110",	-- 105: 	lw	%r1, [%sp + 6]
"00111111111111100000000000000111",	-- 106: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 107: 	addi	%sp, %sp, 8
"01011000000000000010101000011100",	-- 108: 	jal	yj_create_array
"10101011110111100000000000001000",	-- 109: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 110: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000001",	-- 111: 	lli	%r2, 1
"11001100000000110000000000000001",	-- 112: 	lli	%r3, 1
"11001100000001000000000000000000",	-- 113: 	lli	%r4, 0
"10000100001001000010000000000000",	-- 114: 	add	%r4, %r1, %r4
"00111000100001000000000000000000",	-- 115: 	lw	%r4, [%r4 + 0]
"00111100001111100000000000000111",	-- 116: 	sw	%r1, [%sp + 7]
"00111100010111100000000000001000",	-- 117: 	sw	%r2, [%sp + 8]
"10000100000001000001000000000000",	-- 118: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 119: 	add	%r1, %r0, %r3
"00111111111111100000000000001001",	-- 120: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 121: 	addi	%sp, %sp, 10
"01011000000000000010101000011100",	-- 122: 	jal	yj_create_array
"10101011110111100000000000001010",	-- 123: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 124: 	lw	%ra, [%sp + 9]
"10000100000000010001000000000000",	-- 125: 	add	%r2, %r0, %r1
"00111011110000010000000000001000",	-- 126: 	lw	%r1, [%sp + 8]
"00111111111111100000000000001001",	-- 127: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 128: 	addi	%sp, %sp, 10
"01011000000000000010101000011100",	-- 129: 	jal	yj_create_array
"10101011110111100000000000001010",	-- 130: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 131: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000001",	-- 132: 	lli	%r2, 1
"00010100000000000000000000000000",	-- 133: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 134: 	lhif	%f0, 0.000000
"00111100001111100000000000001001",	-- 135: 	sw	%r1, [%sp + 9]
"10000100000000100000100000000000",	-- 136: 	add	%r1, %r0, %r2
"00111111111111100000000000001010",	-- 137: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 138: 	addi	%sp, %sp, 11
"01011000000000000010101000100100",	-- 139: 	jal	yj_create_float_array
"10101011110111100000000000001011",	-- 140: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 141: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000001",	-- 142: 	lli	%r2, 1
"11001100000000110000000000000000",	-- 143: 	lli	%r3, 0
"00111100001111100000000000001010",	-- 144: 	sw	%r1, [%sp + 10]
"10000100000000100000100000000000",	-- 145: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 146: 	add	%r2, %r0, %r3
"00111111111111100000000000001011",	-- 147: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 148: 	addi	%sp, %sp, 12
"01011000000000000010101000011100",	-- 149: 	jal	yj_create_array
"10101011110111100000000000001100",	-- 150: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 151: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000001",	-- 152: 	lli	%r2, 1
"00010100000000000110101100101000",	-- 153: 	llif	%f0, 1000000000.000000
"00010000000000000100111001101110",	-- 154: 	lhif	%f0, 1000000000.000000
"00111100001111100000000000001011",	-- 155: 	sw	%r1, [%sp + 11]
"10000100000000100000100000000000",	-- 156: 	add	%r1, %r0, %r2
"00111111111111100000000000001100",	-- 157: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 158: 	addi	%sp, %sp, 13
"01011000000000000010101000100100",	-- 159: 	jal	yj_create_float_array
"10101011110111100000000000001101",	-- 160: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 161: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000011",	-- 162: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 163: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 164: 	lhif	%f0, 0.000000
"00111100001111100000000000001100",	-- 165: 	sw	%r1, [%sp + 12]
"10000100000000100000100000000000",	-- 166: 	add	%r1, %r0, %r2
"00111111111111100000000000001101",	-- 167: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 168: 	addi	%sp, %sp, 14
"01011000000000000010101000100100",	-- 169: 	jal	yj_create_float_array
"10101011110111100000000000001110",	-- 170: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 171: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000001",	-- 172: 	lli	%r2, 1
"11001100000000110000000000000000",	-- 173: 	lli	%r3, 0
"00111100001111100000000000001101",	-- 174: 	sw	%r1, [%sp + 13]
"10000100000000100000100000000000",	-- 175: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 176: 	add	%r2, %r0, %r3
"00111111111111100000000000001110",	-- 177: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 178: 	addi	%sp, %sp, 15
"01011000000000000010101000011100",	-- 179: 	jal	yj_create_array
"10101011110111100000000000001111",	-- 180: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 181: 	lw	%ra, [%sp + 14]
"11001100000000100000000000000011",	-- 182: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 183: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 184: 	lhif	%f0, 0.000000
"00111100001111100000000000001110",	-- 185: 	sw	%r1, [%sp + 14]
"10000100000000100000100000000000",	-- 186: 	add	%r1, %r0, %r2
"00111111111111100000000000001111",	-- 187: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 188: 	addi	%sp, %sp, 16
"01011000000000000010101000100100",	-- 189: 	jal	yj_create_float_array
"10101011110111100000000000010000",	-- 190: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 191: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000011",	-- 192: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 193: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 194: 	lhif	%f0, 0.000000
"00111100001111100000000000001111",	-- 195: 	sw	%r1, [%sp + 15]
"10000100000000100000100000000000",	-- 196: 	add	%r1, %r0, %r2
"00111111111111100000000000010000",	-- 197: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 198: 	addi	%sp, %sp, 17
"01011000000000000010101000100100",	-- 199: 	jal	yj_create_float_array
"10101011110111100000000000010001",	-- 200: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 201: 	lw	%ra, [%sp + 16]
"11001100000000100000000000000011",	-- 202: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 203: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 204: 	lhif	%f0, 0.000000
"00111100001111100000000000010000",	-- 205: 	sw	%r1, [%sp + 16]
"10000100000000100000100000000000",	-- 206: 	add	%r1, %r0, %r2
"00111111111111100000000000010001",	-- 207: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 208: 	addi	%sp, %sp, 18
"01011000000000000010101000100100",	-- 209: 	jal	yj_create_float_array
"10101011110111100000000000010010",	-- 210: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 211: 	lw	%ra, [%sp + 17]
"11001100000000100000000000000011",	-- 212: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 213: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 214: 	lhif	%f0, 0.000000
"00111100001111100000000000010001",	-- 215: 	sw	%r1, [%sp + 17]
"10000100000000100000100000000000",	-- 216: 	add	%r1, %r0, %r2
"00111111111111100000000000010010",	-- 217: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 218: 	addi	%sp, %sp, 19
"01011000000000000010101000100100",	-- 219: 	jal	yj_create_float_array
"10101011110111100000000000010011",	-- 220: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 221: 	lw	%ra, [%sp + 18]
"11001100000000100000000000000010",	-- 222: 	lli	%r2, 2
"11001100000000110000000000000000",	-- 223: 	lli	%r3, 0
"00111100001111100000000000010010",	-- 224: 	sw	%r1, [%sp + 18]
"10000100000000100000100000000000",	-- 225: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 226: 	add	%r2, %r0, %r3
"00111111111111100000000000010011",	-- 227: 	sw	%ra, [%sp + 19]
"10100111110111100000000000010100",	-- 228: 	addi	%sp, %sp, 20
"01011000000000000010101000011100",	-- 229: 	jal	yj_create_array
"10101011110111100000000000010100",	-- 230: 	subi	%sp, %sp, 20
"00111011110111110000000000010011",	-- 231: 	lw	%ra, [%sp + 19]
"11001100000000100000000000000010",	-- 232: 	lli	%r2, 2
"11001100000000110000000000000000",	-- 233: 	lli	%r3, 0
"00111100001111100000000000010011",	-- 234: 	sw	%r1, [%sp + 19]
"10000100000000100000100000000000",	-- 235: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 236: 	add	%r2, %r0, %r3
"00111111111111100000000000010100",	-- 237: 	sw	%ra, [%sp + 20]
"10100111110111100000000000010101",	-- 238: 	addi	%sp, %sp, 21
"01011000000000000010101000011100",	-- 239: 	jal	yj_create_array
"10101011110111100000000000010101",	-- 240: 	subi	%sp, %sp, 21
"00111011110111110000000000010100",	-- 241: 	lw	%ra, [%sp + 20]
"11001100000000100000000000000001",	-- 242: 	lli	%r2, 1
"00010100000000000000000000000000",	-- 243: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 244: 	lhif	%f0, 0.000000
"00111100001111100000000000010100",	-- 245: 	sw	%r1, [%sp + 20]
"10000100000000100000100000000000",	-- 246: 	add	%r1, %r0, %r2
"00111111111111100000000000010101",	-- 247: 	sw	%ra, [%sp + 21]
"10100111110111100000000000010110",	-- 248: 	addi	%sp, %sp, 22
"01011000000000000010101000100100",	-- 249: 	jal	yj_create_float_array
"10101011110111100000000000010110",	-- 250: 	subi	%sp, %sp, 22
"00111011110111110000000000010101",	-- 251: 	lw	%ra, [%sp + 21]
"11001100000000100000000000000011",	-- 252: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 253: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 254: 	lhif	%f0, 0.000000
"00111100001111100000000000010101",	-- 255: 	sw	%r1, [%sp + 21]
"10000100000000100000100000000000",	-- 256: 	add	%r1, %r0, %r2
"00111111111111100000000000010110",	-- 257: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 258: 	addi	%sp, %sp, 23
"01011000000000000010101000100100",	-- 259: 	jal	yj_create_float_array
"10101011110111100000000000010111",	-- 260: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 261: 	lw	%ra, [%sp + 22]
"11001100000000100000000000000011",	-- 262: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 263: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 264: 	lhif	%f0, 0.000000
"00111100001111100000000000010110",	-- 265: 	sw	%r1, [%sp + 22]
"10000100000000100000100000000000",	-- 266: 	add	%r1, %r0, %r2
"00111111111111100000000000010111",	-- 267: 	sw	%ra, [%sp + 23]
"10100111110111100000000000011000",	-- 268: 	addi	%sp, %sp, 24
"01011000000000000010101000100100",	-- 269: 	jal	yj_create_float_array
"10101011110111100000000000011000",	-- 270: 	subi	%sp, %sp, 24
"00111011110111110000000000010111",	-- 271: 	lw	%ra, [%sp + 23]
"11001100000000100000000000000011",	-- 272: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 273: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 274: 	lhif	%f0, 0.000000
"00111100001111100000000000010111",	-- 275: 	sw	%r1, [%sp + 23]
"10000100000000100000100000000000",	-- 276: 	add	%r1, %r0, %r2
"00111111111111100000000000011000",	-- 277: 	sw	%ra, [%sp + 24]
"10100111110111100000000000011001",	-- 278: 	addi	%sp, %sp, 25
"01011000000000000010101000100100",	-- 279: 	jal	yj_create_float_array
"10101011110111100000000000011001",	-- 280: 	subi	%sp, %sp, 25
"00111011110111110000000000011000",	-- 281: 	lw	%ra, [%sp + 24]
"11001100000000100000000000000011",	-- 282: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 283: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 284: 	lhif	%f0, 0.000000
"00111100001111100000000000011000",	-- 285: 	sw	%r1, [%sp + 24]
"10000100000000100000100000000000",	-- 286: 	add	%r1, %r0, %r2
"00111111111111100000000000011001",	-- 287: 	sw	%ra, [%sp + 25]
"10100111110111100000000000011010",	-- 288: 	addi	%sp, %sp, 26
"01011000000000000010101000100100",	-- 289: 	jal	yj_create_float_array
"10101011110111100000000000011010",	-- 290: 	subi	%sp, %sp, 26
"00111011110111110000000000011001",	-- 291: 	lw	%ra, [%sp + 25]
"11001100000000100000000000000011",	-- 292: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 293: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 294: 	lhif	%f0, 0.000000
"00111100001111100000000000011001",	-- 295: 	sw	%r1, [%sp + 25]
"10000100000000100000100000000000",	-- 296: 	add	%r1, %r0, %r2
"00111111111111100000000000011010",	-- 297: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 298: 	addi	%sp, %sp, 27
"01011000000000000010101000100100",	-- 299: 	jal	yj_create_float_array
"10101011110111100000000000011011",	-- 300: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 301: 	lw	%ra, [%sp + 26]
"11001100000000100000000000000011",	-- 302: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 303: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 304: 	lhif	%f0, 0.000000
"00111100001111100000000000011010",	-- 305: 	sw	%r1, [%sp + 26]
"10000100000000100000100000000000",	-- 306: 	add	%r1, %r0, %r2
"00111111111111100000000000011011",	-- 307: 	sw	%ra, [%sp + 27]
"10100111110111100000000000011100",	-- 308: 	addi	%sp, %sp, 28
"01011000000000000010101000100100",	-- 309: 	jal	yj_create_float_array
"10101011110111100000000000011100",	-- 310: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 311: 	lw	%ra, [%sp + 27]
"11001100000000100000000000000000",	-- 312: 	lli	%r2, 0
"00010100000000000000000000000000",	-- 313: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 314: 	lhif	%f0, 0.000000
"00111100001111100000000000011011",	-- 315: 	sw	%r1, [%sp + 27]
"10000100000000100000100000000000",	-- 316: 	add	%r1, %r0, %r2
"00111111111111100000000000011100",	-- 317: 	sw	%ra, [%sp + 28]
"10100111110111100000000000011101",	-- 318: 	addi	%sp, %sp, 29
"01011000000000000010101000100100",	-- 319: 	jal	yj_create_float_array
"10101011110111100000000000011101",	-- 320: 	subi	%sp, %sp, 29
"00111011110111110000000000011100",	-- 321: 	lw	%ra, [%sp + 28]
"10000100000000010001000000000000",	-- 322: 	add	%r2, %r0, %r1
"11001100000000010000000000000000",	-- 323: 	lli	%r1, 0
"00111100010111100000000000011100",	-- 324: 	sw	%r2, [%sp + 28]
"00111111111111100000000000011101",	-- 325: 	sw	%ra, [%sp + 29]
"10100111110111100000000000011110",	-- 326: 	addi	%sp, %sp, 30
"01011000000000000010101000011100",	-- 327: 	jal	yj_create_array
"10101011110111100000000000011110",	-- 328: 	subi	%sp, %sp, 30
"00111011110111110000000000011101",	-- 329: 	lw	%ra, [%sp + 29]
"11001100000000100000000000000000",	-- 330: 	lli	%r2, 0
"10000100000111010001100000000000",	-- 331: 	add	%r3, %r0, %hp
"10100111101111010000000000000010",	-- 332: 	addi	%hp, %hp, 2
"00111100001000110000000000000001",	-- 333: 	sw	%r1, [%r3 + 1]
"00111011110000010000000000011100",	-- 334: 	lw	%r1, [%sp + 28]
"00111100001000110000000000000000",	-- 335: 	sw	%r1, [%r3 + 0]
"10000100000000110000100000000000",	-- 336: 	add	%r1, %r0, %r3
"10000100000000101101000000000000",	-- 337: 	add	%r26, %r0, %r2
"10000100000000010001000000000000",	-- 338: 	add	%r2, %r0, %r1
"10000100000110100000100000000000",	-- 339: 	add	%r1, %r0, %r26
"00111111111111100000000000011101",	-- 340: 	sw	%ra, [%sp + 29]
"10100111110111100000000000011110",	-- 341: 	addi	%sp, %sp, 30
"01011000000000000010101000011100",	-- 342: 	jal	yj_create_array
"10101011110111100000000000011110",	-- 343: 	subi	%sp, %sp, 30
"00111011110111110000000000011101",	-- 344: 	lw	%ra, [%sp + 29]
"10000100000000010001000000000000",	-- 345: 	add	%r2, %r0, %r1
"11001100000000010000000000000101",	-- 346: 	lli	%r1, 5
"00111111111111100000000000011101",	-- 347: 	sw	%ra, [%sp + 29]
"10100111110111100000000000011110",	-- 348: 	addi	%sp, %sp, 30
"01011000000000000010101000011100",	-- 349: 	jal	yj_create_array
"10101011110111100000000000011110",	-- 350: 	subi	%sp, %sp, 30
"00111011110111110000000000011101",	-- 351: 	lw	%ra, [%sp + 29]
"11001100000000100000000000000000",	-- 352: 	lli	%r2, 0
"00010100000000000000000000000000",	-- 353: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 354: 	lhif	%f0, 0.000000
"00111100001111100000000000011101",	-- 355: 	sw	%r1, [%sp + 29]
"10000100000000100000100000000000",	-- 356: 	add	%r1, %r0, %r2
"00111111111111100000000000011110",	-- 357: 	sw	%ra, [%sp + 30]
"10100111110111100000000000011111",	-- 358: 	addi	%sp, %sp, 31
"01011000000000000010101000100100",	-- 359: 	jal	yj_create_float_array
"10101011110111100000000000011111",	-- 360: 	subi	%sp, %sp, 31
"00111011110111110000000000011110",	-- 361: 	lw	%ra, [%sp + 30]
"11001100000000100000000000000011",	-- 362: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 363: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 364: 	lhif	%f0, 0.000000
"00111100001111100000000000011110",	-- 365: 	sw	%r1, [%sp + 30]
"10000100000000100000100000000000",	-- 366: 	add	%r1, %r0, %r2
"00111111111111100000000000011111",	-- 367: 	sw	%ra, [%sp + 31]
"10100111110111100000000000100000",	-- 368: 	addi	%sp, %sp, 32
"01011000000000000010101000100100",	-- 369: 	jal	yj_create_float_array
"10101011110111100000000000100000",	-- 370: 	subi	%sp, %sp, 32
"00111011110111110000000000011111",	-- 371: 	lw	%ra, [%sp + 31]
"11001100000000100000000000111100",	-- 372: 	lli	%r2, 60
"00111011110000110000000000011110",	-- 373: 	lw	%r3, [%sp + 30]
"00111100001111100000000000011111",	-- 374: 	sw	%r1, [%sp + 31]
"10000100000000100000100000000000",	-- 375: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 376: 	add	%r2, %r0, %r3
"00111111111111100000000000100000",	-- 377: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 378: 	addi	%sp, %sp, 33
"01011000000000000010101000011100",	-- 379: 	jal	yj_create_array
"10101011110111100000000000100001",	-- 380: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 381: 	lw	%ra, [%sp + 32]
"10000100000111010001000000000000",	-- 382: 	add	%r2, %r0, %hp
"10100111101111010000000000000010",	-- 383: 	addi	%hp, %hp, 2
"00111100001000100000000000000001",	-- 384: 	sw	%r1, [%r2 + 1]
"00111011110000010000000000011111",	-- 385: 	lw	%r1, [%sp + 31]
"00111100001000100000000000000000",	-- 386: 	sw	%r1, [%r2 + 0]
"10000100000000100000100000000000",	-- 387: 	add	%r1, %r0, %r2
"11001100000000100000000000000000",	-- 388: 	lli	%r2, 0
"00010100000000000000000000000000",	-- 389: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 390: 	lhif	%f0, 0.000000
"00111100001111100000000000100000",	-- 391: 	sw	%r1, [%sp + 32]
"10000100000000100000100000000000",	-- 392: 	add	%r1, %r0, %r2
"00111111111111100000000000100001",	-- 393: 	sw	%ra, [%sp + 33]
"10100111110111100000000000100010",	-- 394: 	addi	%sp, %sp, 34
"01011000000000000010101000100100",	-- 395: 	jal	yj_create_float_array
"10101011110111100000000000100010",	-- 396: 	subi	%sp, %sp, 34
"00111011110111110000000000100001",	-- 397: 	lw	%ra, [%sp + 33]
"10000100000000010001000000000000",	-- 398: 	add	%r2, %r0, %r1
"11001100000000010000000000000000",	-- 399: 	lli	%r1, 0
"00111100010111100000000000100001",	-- 400: 	sw	%r2, [%sp + 33]
"00111111111111100000000000100010",	-- 401: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 402: 	addi	%sp, %sp, 35
"01011000000000000010101000011100",	-- 403: 	jal	yj_create_array
"10101011110111100000000000100011",	-- 404: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 405: 	lw	%ra, [%sp + 34]
"10000100000111010001000000000000",	-- 406: 	add	%r2, %r0, %hp
"10100111101111010000000000000010",	-- 407: 	addi	%hp, %hp, 2
"00111100001000100000000000000001",	-- 408: 	sw	%r1, [%r2 + 1]
"00111011110000010000000000100001",	-- 409: 	lw	%r1, [%sp + 33]
"00111100001000100000000000000000",	-- 410: 	sw	%r1, [%r2 + 0]
"10000100000000100000100000000000",	-- 411: 	add	%r1, %r0, %r2
"11001100000000100000000010110100",	-- 412: 	lli	%r2, 180
"11001100000000110000000000000000",	-- 413: 	lli	%r3, 0
"00010100000000000000000000000000",	-- 414: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 415: 	lhif	%f0, 0.000000
"10000100000111010010000000000000",	-- 416: 	add	%r4, %r0, %hp
"10100111101111010000000000000011",	-- 417: 	addi	%hp, %hp, 3
"10110000000001000000000000000010",	-- 418: 	sf	%f0, [%r4 + 2]
"00111100001001000000000000000001",	-- 419: 	sw	%r1, [%r4 + 1]
"00111100011001000000000000000000",	-- 420: 	sw	%r3, [%r4 + 0]
"10000100000001000000100000000000",	-- 421: 	add	%r1, %r0, %r4
"10000100000000101101000000000000",	-- 422: 	add	%r26, %r0, %r2
"10000100000000010001000000000000",	-- 423: 	add	%r2, %r0, %r1
"10000100000110100000100000000000",	-- 424: 	add	%r1, %r0, %r26
"00111111111111100000000000100010",	-- 425: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 426: 	addi	%sp, %sp, 35
"01011000000000000010101000011100",	-- 427: 	jal	yj_create_array
"10101011110111100000000000100011",	-- 428: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 429: 	lw	%ra, [%sp + 34]
"11001100000000100000000000000001",	-- 430: 	lli	%r2, 1
"11001100000000110000000000000000",	-- 431: 	lli	%r3, 0
"00111100001111100000000000100010",	-- 432: 	sw	%r1, [%sp + 34]
"10000100000000100000100000000000",	-- 433: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 434: 	add	%r2, %r0, %r3
"00111111111111100000000000100011",	-- 435: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 436: 	addi	%sp, %sp, 36
"01011000000000000010101000011100",	-- 437: 	jal	yj_create_array
"10101011110111100000000000100100",	-- 438: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 439: 	lw	%ra, [%sp + 35]
"10000100000111010001000000000000",	-- 440: 	add	%r2, %r0, %hp
"10100111101111010000000000000110",	-- 441: 	addi	%hp, %hp, 6
"10100100000000110000011011001010",	-- 442: 	addi	%r3, %r0, read_screen_settings.2695
"00111100011000100000000000000000",	-- 443: 	sw	%r3, [%r2 + 0]
"00111011110000110000000000000011",	-- 444: 	lw	%r3, [%sp + 3]
"00111100011000100000000000000101",	-- 445: 	sw	%r3, [%r2 + 5]
"00111011110001000000000000011010",	-- 446: 	lw	%r4, [%sp + 26]
"00111100100000100000000000000100",	-- 447: 	sw	%r4, [%r2 + 4]
"00111011110001010000000000011001",	-- 448: 	lw	%r5, [%sp + 25]
"00111100101000100000000000000011",	-- 449: 	sw	%r5, [%r2 + 3]
"00111011110001100000000000011000",	-- 450: 	lw	%r6, [%sp + 24]
"00111100110000100000000000000010",	-- 451: 	sw	%r6, [%r2 + 2]
"00111011110001110000000000000010",	-- 452: 	lw	%r7, [%sp + 2]
"00111100111000100000000000000001",	-- 453: 	sw	%r7, [%r2 + 1]
"10000100000111010011100000000000",	-- 454: 	add	%r7, %r0, %hp
"10100111101111010000000000000011",	-- 455: 	addi	%hp, %hp, 3
"10100100000010000000011110011101",	-- 456: 	addi	%r8, %r0, read_light.2697
"00111101000001110000000000000000",	-- 457: 	sw	%r8, [%r7 + 0]
"00111011110010000000000000000100",	-- 458: 	lw	%r8, [%sp + 4]
"00111101000001110000000000000010",	-- 459: 	sw	%r8, [%r7 + 2]
"00111011110010010000000000000101",	-- 460: 	lw	%r9, [%sp + 5]
"00111101001001110000000000000001",	-- 461: 	sw	%r9, [%r7 + 1]
"10000100000111010101000000000000",	-- 462: 	add	%r10, %r0, %hp
"10100111101111010000000000000010",	-- 463: 	addi	%hp, %hp, 2
"10100100000010110000100100011100",	-- 464: 	addi	%r11, %r0, read_nth_object.2702
"00111101011010100000000000000000",	-- 465: 	sw	%r11, [%r10 + 0]
"00111011110010110000000000000001",	-- 466: 	lw	%r11, [%sp + 1]
"00111101011010100000000000000001",	-- 467: 	sw	%r11, [%r10 + 1]
"10000100000111010110000000000000",	-- 468: 	add	%r12, %r0, %hp
"10100111101111010000000000000011",	-- 469: 	addi	%hp, %hp, 3
"10100100000011010000101011011001",	-- 470: 	addi	%r13, %r0, read_object.2704
"00111101101011000000000000000000",	-- 471: 	sw	%r13, [%r12 + 0]
"00111101010011000000000000000010",	-- 472: 	sw	%r10, [%r12 + 2]
"00111011110010100000000000000000",	-- 473: 	lw	%r10, [%sp + 0]
"00111101010011000000000000000001",	-- 474: 	sw	%r10, [%r12 + 1]
"10000100000111010110100000000000",	-- 475: 	add	%r13, %r0, %hp
"10100111101111010000000000000010",	-- 476: 	addi	%hp, %hp, 2
"10100100000011100000101011110110",	-- 477: 	addi	%r14, %r0, read_all_object.2706
"00111101110011010000000000000000",	-- 478: 	sw	%r14, [%r13 + 0]
"00111101100011010000000000000001",	-- 479: 	sw	%r12, [%r13 + 1]
"10000100000111010110000000000000",	-- 480: 	add	%r12, %r0, %hp
"10100111101111010000000000000010",	-- 481: 	addi	%hp, %hp, 2
"10100100000011100000101100111001",	-- 482: 	addi	%r14, %r0, read_and_network.2712
"00111101110011000000000000000000",	-- 483: 	sw	%r14, [%r12 + 0]
"00111011110011100000000000000111",	-- 484: 	lw	%r14, [%sp + 7]
"00111101110011000000000000000001",	-- 485: 	sw	%r14, [%r12 + 1]
"10000100000111010111100000000000",	-- 486: 	add	%r15, %r0, %hp
"10100111101111010000000000000110",	-- 487: 	addi	%hp, %hp, 6
"10100100000100000000101101010100",	-- 488: 	addi	%r16, %r0, read_parameter.2714
"00111110000011110000000000000000",	-- 489: 	sw	%r16, [%r15 + 0]
"00111100010011110000000000000101",	-- 490: 	sw	%r2, [%r15 + 5]
"00111100111011110000000000000100",	-- 491: 	sw	%r7, [%r15 + 4]
"00111101100011110000000000000011",	-- 492: 	sw	%r12, [%r15 + 3]
"00111101101011110000000000000010",	-- 493: 	sw	%r13, [%r15 + 2]
"00111011110000100000000000001001",	-- 494: 	lw	%r2, [%sp + 9]
"00111100010011110000000000000001",	-- 495: 	sw	%r2, [%r15 + 1]
"10000100000111010011100000000000",	-- 496: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 497: 	addi	%hp, %hp, 2
"10100100000011000000101110001000",	-- 498: 	addi	%r12, %r0, solver_rect_surface.2716
"00111101100001110000000000000000",	-- 499: 	sw	%r12, [%r7 + 0]
"00111011110011000000000000001010",	-- 500: 	lw	%r12, [%sp + 10]
"00111101100001110000000000000001",	-- 501: 	sw	%r12, [%r7 + 1]
"10000100000111010110100000000000",	-- 502: 	add	%r13, %r0, %hp
"10100111101111010000000000000010",	-- 503: 	addi	%hp, %hp, 2
"10100100000100000000110000001000",	-- 504: 	addi	%r16, %r0, solver_rect.2725
"00111110000011010000000000000000",	-- 505: 	sw	%r16, [%r13 + 0]
"00111100111011010000000000000001",	-- 506: 	sw	%r7, [%r13 + 1]
"10000100000111010011100000000000",	-- 507: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 508: 	addi	%hp, %hp, 2
"10100100000100000000110001000100",	-- 509: 	addi	%r16, %r0, solver_surface.2731
"00111110000001110000000000000000",	-- 510: 	sw	%r16, [%r7 + 0]
"00111101100001110000000000000001",	-- 511: 	sw	%r12, [%r7 + 1]
"10000100000111011000000000000000",	-- 512: 	add	%r16, %r0, %hp
"10100111101111010000000000000010",	-- 513: 	addi	%hp, %hp, 2
"10100100000100010000110101100001",	-- 514: 	addi	%r17, %r0, solver_second.2750
"00111110001100000000000000000000",	-- 515: 	sw	%r17, [%r16 + 0]
"00111101100100000000000000000001",	-- 516: 	sw	%r12, [%r16 + 1]
"10000100000111011000100000000000",	-- 517: 	add	%r17, %r0, %hp
"10100111101111010000000000000101",	-- 518: 	addi	%hp, %hp, 5
"10100100000100100000110111101001",	-- 519: 	addi	%r18, %r0, solver.2756
"00111110010100010000000000000000",	-- 520: 	sw	%r18, [%r17 + 0]
"00111100111100010000000000000100",	-- 521: 	sw	%r7, [%r17 + 4]
"00111110000100010000000000000011",	-- 522: 	sw	%r16, [%r17 + 3]
"00111101101100010000000000000010",	-- 523: 	sw	%r13, [%r17 + 2]
"00111101011100010000000000000001",	-- 524: 	sw	%r11, [%r17 + 1]
"10000100000111010011100000000000",	-- 525: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 526: 	addi	%hp, %hp, 2
"10100100000011010000111000111111",	-- 527: 	addi	%r13, %r0, solver_rect_fast.2760
"00111101101001110000000000000000",	-- 528: 	sw	%r13, [%r7 + 0]
"00111101100001110000000000000001",	-- 529: 	sw	%r12, [%r7 + 1]
"10000100000111010110100000000000",	-- 530: 	add	%r13, %r0, %hp
"10100111101111010000000000000010",	-- 531: 	addi	%hp, %hp, 2
"10100100000100000000111101100101",	-- 532: 	addi	%r16, %r0, solver_surface_fast.2767
"00111110000011010000000000000000",	-- 533: 	sw	%r16, [%r13 + 0]
"00111101100011010000000000000001",	-- 534: 	sw	%r12, [%r13 + 1]
"10000100000111011000000000000000",	-- 535: 	add	%r16, %r0, %hp
"10100111101111010000000000000010",	-- 536: 	addi	%hp, %hp, 2
"10100100000100100000111110010000",	-- 537: 	addi	%r18, %r0, solver_second_fast.2773
"00111110010100000000000000000000",	-- 538: 	sw	%r18, [%r16 + 0]
"00111101100100000000000000000001",	-- 539: 	sw	%r12, [%r16 + 1]
"10000100000111011001000000000000",	-- 540: 	add	%r18, %r0, %hp
"10100111101111010000000000000101",	-- 541: 	addi	%hp, %hp, 5
"10100100000100110001000000010111",	-- 542: 	addi	%r19, %r0, solver_fast.2779
"00111110011100100000000000000000",	-- 543: 	sw	%r19, [%r18 + 0]
"00111101101100100000000000000100",	-- 544: 	sw	%r13, [%r18 + 4]
"00111110000100100000000000000011",	-- 545: 	sw	%r16, [%r18 + 3]
"00111100111100100000000000000010",	-- 546: 	sw	%r7, [%r18 + 2]
"00111101011100100000000000000001",	-- 547: 	sw	%r11, [%r18 + 1]
"10000100000111010110100000000000",	-- 548: 	add	%r13, %r0, %hp
"10100111101111010000000000000010",	-- 549: 	addi	%hp, %hp, 2
"10100100000100000001000010000001",	-- 550: 	addi	%r16, %r0, solver_surface_fast2.2783
"00111110000011010000000000000000",	-- 551: 	sw	%r16, [%r13 + 0]
"00111101100011010000000000000001",	-- 552: 	sw	%r12, [%r13 + 1]
"10000100000111011000000000000000",	-- 553: 	add	%r16, %r0, %hp
"10100111101111010000000000000010",	-- 554: 	addi	%hp, %hp, 2
"10100100000100110001000010100000",	-- 555: 	addi	%r19, %r0, solver_second_fast2.2790
"00111110011100000000000000000000",	-- 556: 	sw	%r19, [%r16 + 0]
"00111101100100000000000000000001",	-- 557: 	sw	%r12, [%r16 + 1]
"10000100000111011001100000000000",	-- 558: 	add	%r19, %r0, %hp
"10100111101111010000000000000101",	-- 559: 	addi	%hp, %hp, 5
"10100100000101000001000100010010",	-- 560: 	addi	%r20, %r0, solver_fast2.2797
"00111110100100110000000000000000",	-- 561: 	sw	%r20, [%r19 + 0]
"00111101101100110000000000000100",	-- 562: 	sw	%r13, [%r19 + 4]
"00111110000100110000000000000011",	-- 563: 	sw	%r16, [%r19 + 3]
"00111100111100110000000000000010",	-- 564: 	sw	%r7, [%r19 + 2]
"00111101011100110000000000000001",	-- 565: 	sw	%r11, [%r19 + 1]
"10000100000111010011100000000000",	-- 566: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 567: 	addi	%hp, %hp, 2
"10100100000011010001001111100011",	-- 568: 	addi	%r13, %r0, iter_setup_dirvec_constants.2809
"00111101101001110000000000000000",	-- 569: 	sw	%r13, [%r7 + 0]
"00111101011001110000000000000001",	-- 570: 	sw	%r11, [%r7 + 1]
"10000100000111010110100000000000",	-- 571: 	add	%r13, %r0, %hp
"10100111101111010000000000000011",	-- 572: 	addi	%hp, %hp, 3
"10100100000100000001010000101111",	-- 573: 	addi	%r16, %r0, setup_dirvec_constants.2812
"00111110000011010000000000000000",	-- 574: 	sw	%r16, [%r13 + 0]
"00111101010011010000000000000010",	-- 575: 	sw	%r10, [%r13 + 2]
"00111100111011010000000000000001",	-- 576: 	sw	%r7, [%r13 + 1]
"10000100000111010011100000000000",	-- 577: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 578: 	addi	%hp, %hp, 2
"10100100000100000001010000111000",	-- 579: 	addi	%r16, %r0, setup_startp_constants.2814
"00111110000001110000000000000000",	-- 580: 	sw	%r16, [%r7 + 0]
"00111101011001110000000000000001",	-- 581: 	sw	%r11, [%r7 + 1]
"10000100000111011000000000000000",	-- 582: 	add	%r16, %r0, %hp
"10100111101111010000000000000100",	-- 583: 	addi	%hp, %hp, 4
"10100100000101000001010011010001",	-- 584: 	addi	%r20, %r0, setup_startp.2817
"00111110100100000000000000000000",	-- 585: 	sw	%r20, [%r16 + 0]
"00111011110101000000000000010111",	-- 586: 	lw	%r20, [%sp + 23]
"00111110100100000000000000000011",	-- 587: 	sw	%r20, [%r16 + 3]
"00111100111100000000000000000010",	-- 588: 	sw	%r7, [%r16 + 2]
"00111101010100000000000000000001",	-- 589: 	sw	%r10, [%r16 + 1]
"10000100000111010011100000000000",	-- 590: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 591: 	addi	%hp, %hp, 2
"10100100000101010001010111010010",	-- 592: 	addi	%r21, %r0, check_all_inside.2839
"00111110101001110000000000000000",	-- 593: 	sw	%r21, [%r7 + 0]
"00111101011001110000000000000001",	-- 594: 	sw	%r11, [%r7 + 1]
"10000100000111011010100000000000",	-- 595: 	add	%r21, %r0, %hp
"10100111101111010000000000001000",	-- 596: 	addi	%hp, %hp, 8
"10100100000101100001010111110110",	-- 597: 	addi	%r22, %r0, shadow_check_and_group.2845
"00111110110101010000000000000000",	-- 598: 	sw	%r22, [%r21 + 0]
"00111110010101010000000000000111",	-- 599: 	sw	%r18, [%r21 + 7]
"00111101100101010000000000000110",	-- 600: 	sw	%r12, [%r21 + 6]
"00111101011101010000000000000101",	-- 601: 	sw	%r11, [%r21 + 5]
"00111011110101100000000000100000",	-- 602: 	lw	%r22, [%sp + 32]
"00111110110101010000000000000100",	-- 603: 	sw	%r22, [%r21 + 4]
"00111101000101010000000000000011",	-- 604: 	sw	%r8, [%r21 + 3]
"00111011110101110000000000001101",	-- 605: 	lw	%r23, [%sp + 13]
"00111110111101010000000000000010",	-- 606: 	sw	%r23, [%r21 + 2]
"00111100111101010000000000000001",	-- 607: 	sw	%r7, [%r21 + 1]
"10000100000111011100000000000000",	-- 608: 	add	%r24, %r0, %hp
"10100111101111010000000000000011",	-- 609: 	addi	%hp, %hp, 3
"10100100000110010001011001110101",	-- 610: 	addi	%r25, %r0, shadow_check_one_or_group.2848
"00111111001110000000000000000000",	-- 611: 	sw	%r25, [%r24 + 0]
"00111110101110000000000000000010",	-- 612: 	sw	%r21, [%r24 + 2]
"00111101110110000000000000000001",	-- 613: 	sw	%r14, [%r24 + 1]
"10000100000111011010100000000000",	-- 614: 	add	%r21, %r0, %hp
"10100111101111010000000000000110",	-- 615: 	addi	%hp, %hp, 6
"10100100000110010001011010011000",	-- 616: 	addi	%r25, %r0, shadow_check_one_or_matrix.2851
"00111111001101010000000000000000",	-- 617: 	sw	%r25, [%r21 + 0]
"00111110010101010000000000000101",	-- 618: 	sw	%r18, [%r21 + 5]
"00111101100101010000000000000100",	-- 619: 	sw	%r12, [%r21 + 4]
"00111111000101010000000000000011",	-- 620: 	sw	%r24, [%r21 + 3]
"00111110110101010000000000000010",	-- 621: 	sw	%r22, [%r21 + 2]
"00111110111101010000000000000001",	-- 622: 	sw	%r23, [%r21 + 1]
"10000100000111011001000000000000",	-- 623: 	add	%r18, %r0, %hp
"10100111101111010000000000001010",	-- 624: 	addi	%hp, %hp, 10
"10100100000110000001011011111001",	-- 625: 	addi	%r24, %r0, solve_each_element.2854
"00111111000100100000000000000000",	-- 626: 	sw	%r24, [%r18 + 0]
"00111011110110000000000000001100",	-- 627: 	lw	%r24, [%sp + 12]
"00111111000100100000000000001001",	-- 628: 	sw	%r24, [%r18 + 9]
"00111011110110010000000000010110",	-- 629: 	lw	%r25, [%sp + 22]
"00111111001100100000000000001000",	-- 630: 	sw	%r25, [%r18 + 8]
"00111101100100100000000000000111",	-- 631: 	sw	%r12, [%r18 + 7]
"00111110001100100000000000000110",	-- 632: 	sw	%r17, [%r18 + 6]
"00111101011100100000000000000101",	-- 633: 	sw	%r11, [%r18 + 5]
"00111011110110100000000000001011",	-- 634: 	lw	%r26, [%sp + 11]
"00111111010100100000000000000100",	-- 635: 	sw	%r26, [%r18 + 4]
"00111110111100100000000000000011",	-- 636: 	sw	%r23, [%r18 + 3]
"00111011110110110000000000001110",	-- 637: 	lw	%r27, [%sp + 14]
"00111111011100100000000000000010",	-- 638: 	sw	%r27, [%r18 + 2]
"00111100111100100000000000000001",	-- 639: 	sw	%r7, [%r18 + 1]
"10000100000111011011000000000000",	-- 640: 	add	%r22, %r0, %hp
"10100111101111010000000000000011",	-- 641: 	addi	%hp, %hp, 3
"00111101111111100000000000100011",	-- 642: 	sw	%r15, [%sp + 35]
"10100100000011110001011110100100",	-- 643: 	addi	%r15, %r0, solve_one_or_network.2858
"00111101111101100000000000000000",	-- 644: 	sw	%r15, [%r22 + 0]
"00111110010101100000000000000010",	-- 645: 	sw	%r18, [%r22 + 2]
"00111101110101100000000000000001",	-- 646: 	sw	%r14, [%r22 + 1]
"10000100000111010111100000000000",	-- 647: 	add	%r15, %r0, %hp
"10100111101111010000000000000110",	-- 648: 	addi	%hp, %hp, 6
"10100100000100100001011111000100",	-- 649: 	addi	%r18, %r0, trace_or_matrix.2862
"00111110010011110000000000000000",	-- 650: 	sw	%r18, [%r15 + 0]
"00111111000011110000000000000101",	-- 651: 	sw	%r24, [%r15 + 5]
"00111111001011110000000000000100",	-- 652: 	sw	%r25, [%r15 + 4]
"00111101100011110000000000000011",	-- 653: 	sw	%r12, [%r15 + 3]
"00111110001011110000000000000010",	-- 654: 	sw	%r17, [%r15 + 2]
"00111110110011110000000000000001",	-- 655: 	sw	%r22, [%r15 + 1]
"10000100000111011000100000000000",	-- 656: 	add	%r17, %r0, %hp
"10100111101111010000000000000100",	-- 657: 	addi	%hp, %hp, 4
"10100100000100100001100000010110",	-- 658: 	addi	%r18, %r0, judge_intersection.2866
"00111110010100010000000000000000",	-- 659: 	sw	%r18, [%r17 + 0]
"00111101111100010000000000000011",	-- 660: 	sw	%r15, [%r17 + 3]
"00111111000100010000000000000010",	-- 661: 	sw	%r24, [%r17 + 2]
"00111100010100010000000000000001",	-- 662: 	sw	%r2, [%r17 + 1]
"10000100000111010111100000000000",	-- 663: 	add	%r15, %r0, %hp
"10100111101111010000000000001010",	-- 664: 	addi	%hp, %hp, 10
"10100100000100100001100001000001",	-- 665: 	addi	%r18, %r0, solve_each_element_fast.2868
"00111110010011110000000000000000",	-- 666: 	sw	%r18, [%r15 + 0]
"00111111000011110000000000001001",	-- 667: 	sw	%r24, [%r15 + 9]
"00111110100011110000000000001000",	-- 668: 	sw	%r20, [%r15 + 8]
"00111110011011110000000000000111",	-- 669: 	sw	%r19, [%r15 + 7]
"00111101100011110000000000000110",	-- 670: 	sw	%r12, [%r15 + 6]
"00111101011011110000000000000101",	-- 671: 	sw	%r11, [%r15 + 5]
"00111111010011110000000000000100",	-- 672: 	sw	%r26, [%r15 + 4]
"00111110111011110000000000000011",	-- 673: 	sw	%r23, [%r15 + 3]
"00111111011011110000000000000010",	-- 674: 	sw	%r27, [%r15 + 2]
"00111100111011110000000000000001",	-- 675: 	sw	%r7, [%r15 + 1]
"10000100000111010011100000000000",	-- 676: 	add	%r7, %r0, %hp
"10100111101111010000000000000011",	-- 677: 	addi	%hp, %hp, 3
"10100100000100100001100011110101",	-- 678: 	addi	%r18, %r0, solve_one_or_network_fast.2872
"00111110010001110000000000000000",	-- 679: 	sw	%r18, [%r7 + 0]
"00111101111001110000000000000010",	-- 680: 	sw	%r15, [%r7 + 2]
"00111101110001110000000000000001",	-- 681: 	sw	%r14, [%r7 + 1]
"10000100000111010111000000000000",	-- 682: 	add	%r14, %r0, %hp
"10100111101111010000000000000101",	-- 683: 	addi	%hp, %hp, 5
"10100100000011110001100100010101",	-- 684: 	addi	%r15, %r0, trace_or_matrix_fast.2876
"00111101111011100000000000000000",	-- 685: 	sw	%r15, [%r14 + 0]
"00111111000011100000000000000100",	-- 686: 	sw	%r24, [%r14 + 4]
"00111110011011100000000000000011",	-- 687: 	sw	%r19, [%r14 + 3]
"00111101100011100000000000000010",	-- 688: 	sw	%r12, [%r14 + 2]
"00111100111011100000000000000001",	-- 689: 	sw	%r7, [%r14 + 1]
"10000100000111010011100000000000",	-- 690: 	add	%r7, %r0, %hp
"10100111101111010000000000000100",	-- 691: 	addi	%hp, %hp, 4
"10100100000011000001100101100101",	-- 692: 	addi	%r12, %r0, judge_intersection_fast.2880
"00111101100001110000000000000000",	-- 693: 	sw	%r12, [%r7 + 0]
"00111101110001110000000000000011",	-- 694: 	sw	%r14, [%r7 + 3]
"00111111000001110000000000000010",	-- 695: 	sw	%r24, [%r7 + 2]
"00111100010001110000000000000001",	-- 696: 	sw	%r2, [%r7 + 1]
"10000100000111010110000000000000",	-- 697: 	add	%r12, %r0, %hp
"10100111101111010000000000000011",	-- 698: 	addi	%hp, %hp, 3
"10100100000011100001100110010000",	-- 699: 	addi	%r14, %r0, get_nvector_rect.2882
"00111101110011000000000000000000",	-- 700: 	sw	%r14, [%r12 + 0]
"00111011110011100000000000001111",	-- 701: 	lw	%r14, [%sp + 15]
"00111101110011000000000000000010",	-- 702: 	sw	%r14, [%r12 + 2]
"00111111010011000000000000000001",	-- 703: 	sw	%r26, [%r12 + 1]
"10000100000111010111100000000000",	-- 704: 	add	%r15, %r0, %hp
"10100111101111010000000000000010",	-- 705: 	addi	%hp, %hp, 2
"10100100000100100001100110110110",	-- 706: 	addi	%r18, %r0, get_nvector_plane.2884
"00111110010011110000000000000000",	-- 707: 	sw	%r18, [%r15 + 0]
"00111101110011110000000000000001",	-- 708: 	sw	%r14, [%r15 + 1]
"10000100000111011001000000000000",	-- 709: 	add	%r18, %r0, %hp
"10100111101111010000000000000011",	-- 710: 	addi	%hp, %hp, 3
"10100100000100110001100111101110",	-- 711: 	addi	%r19, %r0, get_nvector_second.2886
"00111110011100100000000000000000",	-- 712: 	sw	%r19, [%r18 + 0]
"00111101110100100000000000000010",	-- 713: 	sw	%r14, [%r18 + 2]
"00111110111100100000000000000001",	-- 714: 	sw	%r23, [%r18 + 1]
"10000100000111011001100000000000",	-- 715: 	add	%r19, %r0, %hp
"10100111101111010000000000000100",	-- 716: 	addi	%hp, %hp, 4
"10100100000101000001101010111000",	-- 717: 	addi	%r20, %r0, get_nvector.2888
"00111110100100110000000000000000",	-- 718: 	sw	%r20, [%r19 + 0]
"00111110010100110000000000000011",	-- 719: 	sw	%r18, [%r19 + 3]
"00111101100100110000000000000010",	-- 720: 	sw	%r12, [%r19 + 2]
"00111101111100110000000000000001",	-- 721: 	sw	%r15, [%r19 + 1]
"10000100000111010110000000000000",	-- 722: 	add	%r12, %r0, %hp
"10100111101111010000000000000010",	-- 723: 	addi	%hp, %hp, 2
"10100100000011110001101011010101",	-- 724: 	addi	%r15, %r0, utexture.2891
"00111101111011000000000000000000",	-- 725: 	sw	%r15, [%r12 + 0]
"00111011110011110000000000010000",	-- 726: 	lw	%r15, [%sp + 16]
"00111101111011000000000000000001",	-- 727: 	sw	%r15, [%r12 + 1]
"10000100000111011001000000000000",	-- 728: 	add	%r18, %r0, %hp
"10100111101111010000000000000011",	-- 729: 	addi	%hp, %hp, 3
"10100100000101000001110011100011",	-- 730: 	addi	%r20, %r0, add_light.2894
"00111110100100100000000000000000",	-- 731: 	sw	%r20, [%r18 + 0]
"00111101111100100000000000000010",	-- 732: 	sw	%r15, [%r18 + 2]
"00111011110101000000000000010010",	-- 733: 	lw	%r20, [%sp + 18]
"00111110100100100000000000000001",	-- 734: 	sw	%r20, [%r18 + 1]
"10000100000111011011000000000000",	-- 735: 	add	%r22, %r0, %hp
"10100111101111010000000000001001",	-- 736: 	addi	%hp, %hp, 9
"00111101101111100000000000100100",	-- 737: 	sw	%r13, [%sp + 36]
"10100100000011010001110100100111",	-- 738: 	addi	%r13, %r0, trace_reflections.2898
"00111101101101100000000000000000",	-- 739: 	sw	%r13, [%r22 + 0]
"00111110101101100000000000001000",	-- 740: 	sw	%r21, [%r22 + 8]
"00111011110011010000000000100010",	-- 741: 	lw	%r13, [%sp + 34]
"00111101101101100000000000000111",	-- 742: 	sw	%r13, [%r22 + 7]
"00111100010101100000000000000110",	-- 743: 	sw	%r2, [%r22 + 6]
"00111101110101100000000000000101",	-- 744: 	sw	%r14, [%r22 + 5]
"00111100111101100000000000000100",	-- 745: 	sw	%r7, [%r22 + 4]
"00111111010101100000000000000011",	-- 746: 	sw	%r26, [%r22 + 3]
"00111111011101100000000000000010",	-- 747: 	sw	%r27, [%r22 + 2]
"00111110010101100000000000000001",	-- 748: 	sw	%r18, [%r22 + 1]
"10000100000111010110100000000000",	-- 749: 	add	%r13, %r0, %hp
"10100111101111010000000000010101",	-- 750: 	addi	%hp, %hp, 21
"10100100000010100001110110110010",	-- 751: 	addi	%r10, %r0, trace_ray.2903
"00111101010011010000000000000000",	-- 752: 	sw	%r10, [%r13 + 0]
"00111101100011010000000000010100",	-- 753: 	sw	%r12, [%r13 + 20]
"00111110110011010000000000010011",	-- 754: 	sw	%r22, [%r13 + 19]
"00111111000011010000000000010010",	-- 755: 	sw	%r24, [%r13 + 18]
"00111101111011010000000000010001",	-- 756: 	sw	%r15, [%r13 + 17]
"00111111001011010000000000010000",	-- 757: 	sw	%r25, [%r13 + 16]
"00111110101011010000000000001111",	-- 758: 	sw	%r21, [%r13 + 15]
"00111110000011010000000000001110",	-- 759: 	sw	%r16, [%r13 + 14]
"00111110100011010000000000001101",	-- 760: 	sw	%r20, [%r13 + 13]
"00111100010011010000000000001100",	-- 761: 	sw	%r2, [%r13 + 12]
"00111101011011010000000000001011",	-- 762: 	sw	%r11, [%r13 + 11]
"00111101110011010000000000001010",	-- 763: 	sw	%r14, [%r13 + 10]
"00111100001011010000000000001001",	-- 764: 	sw	%r1, [%r13 + 9]
"00111101000011010000000000001000",	-- 765: 	sw	%r8, [%r13 + 8]
"00111110001011010000000000000111",	-- 766: 	sw	%r17, [%r13 + 7]
"00111111010011010000000000000110",	-- 767: 	sw	%r26, [%r13 + 6]
"00111110111011010000000000000101",	-- 768: 	sw	%r23, [%r13 + 5]
"00111111011011010000000000000100",	-- 769: 	sw	%r27, [%r13 + 4]
"00111110011011010000000000000011",	-- 770: 	sw	%r19, [%r13 + 3]
"00111101001011010000000000000010",	-- 771: 	sw	%r9, [%r13 + 2]
"00111110010011010000000000000001",	-- 772: 	sw	%r18, [%r13 + 1]
"10000100000111010100100000000000",	-- 773: 	add	%r9, %r0, %hp
"10100111101111010000000000001101",	-- 774: 	addi	%hp, %hp, 13
"10100100000010100001111101110111",	-- 775: 	addi	%r10, %r0, trace_diffuse_ray.2909
"00111101010010010000000000000000",	-- 776: 	sw	%r10, [%r9 + 0]
"00111101100010010000000000001100",	-- 777: 	sw	%r12, [%r9 + 12]
"00111101111010010000000000001011",	-- 778: 	sw	%r15, [%r9 + 11]
"00111110101010010000000000001010",	-- 779: 	sw	%r21, [%r9 + 10]
"00111100010010010000000000001001",	-- 780: 	sw	%r2, [%r9 + 9]
"00111101011010010000000000001000",	-- 781: 	sw	%r11, [%r9 + 8]
"00111101110010010000000000000111",	-- 782: 	sw	%r14, [%r9 + 7]
"00111101000010010000000000000110",	-- 783: 	sw	%r8, [%r9 + 6]
"00111100111010010000000000000101",	-- 784: 	sw	%r7, [%r9 + 5]
"00111110111010010000000000000100",	-- 785: 	sw	%r23, [%r9 + 4]
"00111111011010010000000000000011",	-- 786: 	sw	%r27, [%r9 + 3]
"00111110011010010000000000000010",	-- 787: 	sw	%r19, [%r9 + 2]
"00111011110000100000000000010001",	-- 788: 	lw	%r2, [%sp + 17]
"00111100010010010000000000000001",	-- 789: 	sw	%r2, [%r9 + 1]
"10000100000111010011100000000000",	-- 790: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 791: 	addi	%hp, %hp, 2
"10100100000010100001111111110000",	-- 792: 	addi	%r10, %r0, iter_trace_diffuse_rays.2912
"00111101010001110000000000000000",	-- 793: 	sw	%r10, [%r7 + 0]
"00111101001001110000000000000001",	-- 794: 	sw	%r9, [%r7 + 1]
"10000100000111010100100000000000",	-- 795: 	add	%r9, %r0, %hp
"10100111101111010000000000000011",	-- 796: 	addi	%hp, %hp, 3
"10100100000010100010000000111011",	-- 797: 	addi	%r10, %r0, trace_diffuse_rays.2917
"00111101010010010000000000000000",	-- 798: 	sw	%r10, [%r9 + 0]
"00111110000010010000000000000010",	-- 799: 	sw	%r16, [%r9 + 2]
"00111100111010010000000000000001",	-- 800: 	sw	%r7, [%r9 + 1]
"10000100000111010011100000000000",	-- 801: 	add	%r7, %r0, %hp
"10100111101111010000000000000011",	-- 802: 	addi	%hp, %hp, 3
"10100100000010100010000001010000",	-- 803: 	addi	%r10, %r0, trace_diffuse_ray_80percent.2921
"00111101010001110000000000000000",	-- 804: 	sw	%r10, [%r7 + 0]
"00111101001001110000000000000010",	-- 805: 	sw	%r9, [%r7 + 2]
"00111011110010100000000000011101",	-- 806: 	lw	%r10, [%sp + 29]
"00111101010001110000000000000001",	-- 807: 	sw	%r10, [%r7 + 1]
"10000100000111010110000000000000",	-- 808: 	add	%r12, %r0, %hp
"10100111101111010000000000000100",	-- 809: 	addi	%hp, %hp, 4
"10100100000011100010000010101011",	-- 810: 	addi	%r14, %r0, calc_diffuse_using_1point.2925
"00111101110011000000000000000000",	-- 811: 	sw	%r14, [%r12 + 0]
"00111100111011000000000000000011",	-- 812: 	sw	%r7, [%r12 + 3]
"00111110100011000000000000000010",	-- 813: 	sw	%r20, [%r12 + 2]
"00111100010011000000000000000001",	-- 814: 	sw	%r2, [%r12 + 1]
"10000100000111010011100000000000",	-- 815: 	add	%r7, %r0, %hp
"10100111101111010000000000000011",	-- 816: 	addi	%hp, %hp, 3
"10100100000011100010000011111010",	-- 817: 	addi	%r14, %r0, calc_diffuse_using_5points.2928
"00111101110001110000000000000000",	-- 818: 	sw	%r14, [%r7 + 0]
"00111110100001110000000000000010",	-- 819: 	sw	%r20, [%r7 + 2]
"00111100010001110000000000000001",	-- 820: 	sw	%r2, [%r7 + 1]
"10000100000111010111000000000000",	-- 821: 	add	%r14, %r0, %hp
"10100111101111010000000000000010",	-- 822: 	addi	%hp, %hp, 2
"10100100000011110010000110000010",	-- 823: 	addi	%r15, %r0, do_without_neighbors.2934
"00111101111011100000000000000000",	-- 824: 	sw	%r15, [%r14 + 0]
"00111101100011100000000000000001",	-- 825: 	sw	%r12, [%r14 + 1]
"10000100000111010110000000000000",	-- 826: 	add	%r12, %r0, %hp
"10100111101111010000000000000010",	-- 827: 	addi	%hp, %hp, 2
"10100100000011110010000110110000",	-- 828: 	addi	%r15, %r0, neighbors_exist.2937
"00111101111011000000000000000000",	-- 829: 	sw	%r15, [%r12 + 0]
"00111011110011110000000000010011",	-- 830: 	lw	%r15, [%sp + 19]
"00111101111011000000000000000001",	-- 831: 	sw	%r15, [%r12 + 1]
"10000100000111011000000000000000",	-- 832: 	add	%r16, %r0, %hp
"10100111101111010000000000000011",	-- 833: 	addi	%hp, %hp, 3
"10100100000100010010001000101000",	-- 834: 	addi	%r17, %r0, try_exploit_neighbors.2950
"00111110001100000000000000000000",	-- 835: 	sw	%r17, [%r16 + 0]
"00111101110100000000000000000010",	-- 836: 	sw	%r14, [%r16 + 2]
"00111100111100000000000000000001",	-- 837: 	sw	%r7, [%r16 + 1]
"10000100000111010011100000000000",	-- 838: 	add	%r7, %r0, %hp
"10100111101111010000000000000010",	-- 839: 	addi	%hp, %hp, 2
"10100100000100010010001001111011",	-- 840: 	addi	%r17, %r0, write_ppm_header.2957
"00111110001001110000000000000000",	-- 841: 	sw	%r17, [%r7 + 0]
"00111101111001110000000000000001",	-- 842: 	sw	%r15, [%r7 + 1]
"10000100000111011000100000000000",	-- 843: 	add	%r17, %r0, %hp
"10100111101111010000000000000010",	-- 844: 	addi	%hp, %hp, 2
"10100100000100100010001011000100",	-- 845: 	addi	%r18, %r0, write_rgb.2961
"00111110010100010000000000000000",	-- 846: 	sw	%r18, [%r17 + 0]
"00111110100100010000000000000001",	-- 847: 	sw	%r20, [%r17 + 1]
"10000100000111011001000000000000",	-- 848: 	add	%r18, %r0, %hp
"10100111101111010000000000000100",	-- 849: 	addi	%hp, %hp, 4
"10100100000100110010001011101110",	-- 850: 	addi	%r19, %r0, pretrace_diffuse_rays.2963
"00111110011100100000000000000000",	-- 851: 	sw	%r19, [%r18 + 0]
"00111101001100100000000000000011",	-- 852: 	sw	%r9, [%r18 + 3]
"00111101010100100000000000000010",	-- 853: 	sw	%r10, [%r18 + 2]
"00111100010100100000000000000001",	-- 854: 	sw	%r2, [%r18 + 1]
"10000100000111010001000000000000",	-- 855: 	add	%r2, %r0, %hp
"10100111101111010000000000001010",	-- 856: 	addi	%hp, %hp, 10
"10100100000010010010001101010101",	-- 857: 	addi	%r9, %r0, pretrace_pixels.2966
"00111101001000100000000000000000",	-- 858: 	sw	%r9, [%r2 + 0]
"00111100011000100000000000001001",	-- 859: 	sw	%r3, [%r2 + 9]
"00111101101000100000000000001000",	-- 860: 	sw	%r13, [%r2 + 8]
"00111111001000100000000000000111",	-- 861: 	sw	%r25, [%r2 + 7]
"00111100110000100000000000000110",	-- 862: 	sw	%r6, [%r2 + 6]
"00111011110000110000000000010101",	-- 863: 	lw	%r3, [%sp + 21]
"00111100011000100000000000000101",	-- 864: 	sw	%r3, [%r2 + 5]
"00111110100000100000000000000100",	-- 865: 	sw	%r20, [%r2 + 4]
"00111011110001100000000000011011",	-- 866: 	lw	%r6, [%sp + 27]
"00111100110000100000000000000011",	-- 867: 	sw	%r6, [%r2 + 3]
"00111110010000100000000000000010",	-- 868: 	sw	%r18, [%r2 + 2]
"00111011110001100000000000010100",	-- 869: 	lw	%r6, [%sp + 20]
"00111100110000100000000000000001",	-- 870: 	sw	%r6, [%r2 + 1]
"10000100000111010100100000000000",	-- 871: 	add	%r9, %r0, %hp
"10100111101111010000000000000111",	-- 872: 	addi	%hp, %hp, 7
"10100100000011010010010000000100",	-- 873: 	addi	%r13, %r0, pretrace_line.2973
"00111101101010010000000000000000",	-- 874: 	sw	%r13, [%r9 + 0]
"00111100100010010000000000000110",	-- 875: 	sw	%r4, [%r9 + 6]
"00111100101010010000000000000101",	-- 876: 	sw	%r5, [%r9 + 5]
"00111100011010010000000000000100",	-- 877: 	sw	%r3, [%r9 + 4]
"00111100010010010000000000000011",	-- 878: 	sw	%r2, [%r9 + 3]
"00111101111010010000000000000010",	-- 879: 	sw	%r15, [%r9 + 2]
"00111100110010010000000000000001",	-- 880: 	sw	%r6, [%r9 + 1]
"10000100000111010001000000000000",	-- 881: 	add	%r2, %r0, %hp
"10100111101111010000000000000111",	-- 882: 	addi	%hp, %hp, 7
"10100100000001000010010001001001",	-- 883: 	addi	%r4, %r0, scan_pixel.2977
"00111100100000100000000000000000",	-- 884: 	sw	%r4, [%r2 + 0]
"00111110001000100000000000000110",	-- 885: 	sw	%r17, [%r2 + 6]
"00111110000000100000000000000101",	-- 886: 	sw	%r16, [%r2 + 5]
"00111110100000100000000000000100",	-- 887: 	sw	%r20, [%r2 + 4]
"00111101100000100000000000000011",	-- 888: 	sw	%r12, [%r2 + 3]
"00111101111000100000000000000010",	-- 889: 	sw	%r15, [%r2 + 2]
"00111101110000100000000000000001",	-- 890: 	sw	%r14, [%r2 + 1]
"10000100000111010010000000000000",	-- 891: 	add	%r4, %r0, %hp
"10100111101111010000000000000100",	-- 892: 	addi	%hp, %hp, 4
"10100100000001010010010010100111",	-- 893: 	addi	%r5, %r0, scan_line.2983
"00111100101001000000000000000000",	-- 894: 	sw	%r5, [%r4 + 0]
"00111100010001000000000000000011",	-- 895: 	sw	%r2, [%r4 + 3]
"00111101001001000000000000000010",	-- 896: 	sw	%r9, [%r4 + 2]
"00111101111001000000000000000001",	-- 897: 	sw	%r15, [%r4 + 1]
"10000100000111010001000000000000",	-- 898: 	add	%r2, %r0, %hp
"10100111101111010000000000000010",	-- 899: 	addi	%hp, %hp, 2
"10100100000001010010010110011010",	-- 900: 	addi	%r5, %r0, create_pixelline.2996
"00111100101000100000000000000000",	-- 901: 	sw	%r5, [%r2 + 0]
"00111101111000100000000000000001",	-- 902: 	sw	%r15, [%r2 + 1]
"10000100000111010010100000000000",	-- 903: 	add	%r5, %r0, %hp
"10100111101111010000000000000010",	-- 904: 	addi	%hp, %hp, 2
"10100100000011000010010111100010",	-- 905: 	addi	%r12, %r0, calc_dirvec.3003
"00111101100001010000000000000000",	-- 906: 	sw	%r12, [%r5 + 0]
"00111101010001010000000000000001",	-- 907: 	sw	%r10, [%r5 + 1]
"10000100000111010110000000000000",	-- 908: 	add	%r12, %r0, %hp
"10100111101111010000000000000010",	-- 909: 	addi	%hp, %hp, 2
"10100100000011010010011011100101",	-- 910: 	addi	%r13, %r0, calc_dirvecs.3011
"00111101101011000000000000000000",	-- 911: 	sw	%r13, [%r12 + 0]
"00111100101011000000000000000001",	-- 912: 	sw	%r5, [%r12 + 1]
"10000100000111010010100000000000",	-- 913: 	add	%r5, %r0, %hp
"10100111101111010000000000000010",	-- 914: 	addi	%hp, %hp, 2
"10100100000011010010011100111011",	-- 915: 	addi	%r13, %r0, calc_dirvec_rows.3016
"00111101101001010000000000000000",	-- 916: 	sw	%r13, [%r5 + 0]
"00111101100001010000000000000001",	-- 917: 	sw	%r12, [%r5 + 1]
"10000100000111010110000000000000",	-- 918: 	add	%r12, %r0, %hp
"10100111101111010000000000000010",	-- 919: 	addi	%hp, %hp, 2
"10100100000011010010011101101101",	-- 920: 	addi	%r13, %r0, create_dirvec.3020
"00111101101011000000000000000000",	-- 921: 	sw	%r13, [%r12 + 0]
"00111011110011010000000000000000",	-- 922: 	lw	%r13, [%sp + 0]
"00111101101011000000000000000001",	-- 923: 	sw	%r13, [%r12 + 1]
"10000100000111010111000000000000",	-- 924: 	add	%r14, %r0, %hp
"10100111101111010000000000000010",	-- 925: 	addi	%hp, %hp, 2
"10100100000100000010011110001010",	-- 926: 	addi	%r16, %r0, create_dirvec_elements.3022
"00111110000011100000000000000000",	-- 927: 	sw	%r16, [%r14 + 0]
"00111101100011100000000000000001",	-- 928: 	sw	%r12, [%r14 + 1]
"10000100000111011000000000000000",	-- 929: 	add	%r16, %r0, %hp
"10100111101111010000000000000100",	-- 930: 	addi	%hp, %hp, 4
"10100100000100010010011110100010",	-- 931: 	addi	%r17, %r0, create_dirvecs.3025
"00111110001100000000000000000000",	-- 932: 	sw	%r17, [%r16 + 0]
"00111101010100000000000000000011",	-- 933: 	sw	%r10, [%r16 + 3]
"00111101110100000000000000000010",	-- 934: 	sw	%r14, [%r16 + 2]
"00111101100100000000000000000001",	-- 935: 	sw	%r12, [%r16 + 1]
"10000100000111010111000000000000",	-- 936: 	add	%r14, %r0, %hp
"10100111101111010000000000000010",	-- 937: 	addi	%hp, %hp, 2
"10100100000100010010011111010001",	-- 938: 	addi	%r17, %r0, init_dirvec_constants.3027
"00111110001011100000000000000000",	-- 939: 	sw	%r17, [%r14 + 0]
"00111011110100010000000000100100",	-- 940: 	lw	%r17, [%sp + 36]
"00111110001011100000000000000001",	-- 941: 	sw	%r17, [%r14 + 1]
"10000100000111011001000000000000",	-- 942: 	add	%r18, %r0, %hp
"10100111101111010000000000000011",	-- 943: 	addi	%hp, %hp, 3
"10100100000100110010011111101001",	-- 944: 	addi	%r19, %r0, init_vecset_constants.3030
"00111110011100100000000000000000",	-- 945: 	sw	%r19, [%r18 + 0]
"00111101110100100000000000000010",	-- 946: 	sw	%r14, [%r18 + 2]
"00111101010100100000000000000001",	-- 947: 	sw	%r10, [%r18 + 1]
"10000100000111010101000000000000",	-- 948: 	add	%r10, %r0, %hp
"10100111101111010000000000000100",	-- 949: 	addi	%hp, %hp, 4
"10100100000011100010100000000010",	-- 950: 	addi	%r14, %r0, init_dirvecs.3032
"00111101110010100000000000000000",	-- 951: 	sw	%r14, [%r10 + 0]
"00111110010010100000000000000011",	-- 952: 	sw	%r18, [%r10 + 3]
"00111110000010100000000000000010",	-- 953: 	sw	%r16, [%r10 + 2]
"00111100101010100000000000000001",	-- 954: 	sw	%r5, [%r10 + 1]
"10000100000111010010100000000000",	-- 955: 	add	%r5, %r0, %hp
"10100111101111010000000000000100",	-- 956: 	addi	%hp, %hp, 4
"10100100000011100010100000011110",	-- 957: 	addi	%r14, %r0, add_reflection.3034
"00111101110001010000000000000000",	-- 958: 	sw	%r14, [%r5 + 0]
"00111110001001010000000000000011",	-- 959: 	sw	%r17, [%r5 + 3]
"00111011110011100000000000100010",	-- 960: 	lw	%r14, [%sp + 34]
"00111101110001010000000000000010",	-- 961: 	sw	%r14, [%r5 + 2]
"00111101100001010000000000000001",	-- 962: 	sw	%r12, [%r5 + 1]
"10000100000111010110000000000000",	-- 963: 	add	%r12, %r0, %hp
"10100111101111010000000000000100",	-- 964: 	addi	%hp, %hp, 4
"10100100000011100010100001010010",	-- 965: 	addi	%r14, %r0, setup_rect_reflection.3041
"00111101110011000000000000000000",	-- 966: 	sw	%r14, [%r12 + 0]
"00111100001011000000000000000011",	-- 967: 	sw	%r1, [%r12 + 3]
"00111101000011000000000000000010",	-- 968: 	sw	%r8, [%r12 + 2]
"00111100101011000000000000000001",	-- 969: 	sw	%r5, [%r12 + 1]
"10000100000111010111000000000000",	-- 970: 	add	%r14, %r0, %hp
"10100111101111010000000000000100",	-- 971: 	addi	%hp, %hp, 4
"10100100000100000010100011010010",	-- 972: 	addi	%r16, %r0, setup_surface_reflection.3044
"00111110000011100000000000000000",	-- 973: 	sw	%r16, [%r14 + 0]
"00111100001011100000000000000011",	-- 974: 	sw	%r1, [%r14 + 3]
"00111101000011100000000000000010",	-- 975: 	sw	%r8, [%r14 + 2]
"00111100101011100000000000000001",	-- 976: 	sw	%r5, [%r14 + 1]
"10000100000111010000100000000000",	-- 977: 	add	%r1, %r0, %hp
"10100111101111010000000000000100",	-- 978: 	addi	%hp, %hp, 4
"10100100000001010010100101001000",	-- 979: 	addi	%r5, %r0, setup_reflections.3047
"00111100101000010000000000000000",	-- 980: 	sw	%r5, [%r1 + 0]
"00111101110000010000000000000011",	-- 981: 	sw	%r14, [%r1 + 3]
"00111101100000010000000000000010",	-- 982: 	sw	%r12, [%r1 + 2]
"00111101011000010000000000000001",	-- 983: 	sw	%r11, [%r1 + 1]
"10000100000111011101100000000000",	-- 984: 	add	%r27, %r0, %hp
"10100111101111010000000000001111",	-- 985: 	addi	%hp, %hp, 15
"10100100000001010010100110000010",	-- 986: 	addi	%r5, %r0, rt.3049
"00111100101110110000000000000000",	-- 987: 	sw	%r5, [%r27 + 0]
"00111100111110110000000000001110",	-- 988: 	sw	%r7, [%r27 + 14]
"00111100001110110000000000001101",	-- 989: 	sw	%r1, [%r27 + 13]
"00111110001110110000000000001100",	-- 990: 	sw	%r17, [%r27 + 12]
"00111100011110110000000000001011",	-- 991: 	sw	%r3, [%r27 + 11]
"00111100100110110000000000001010",	-- 992: 	sw	%r4, [%r27 + 10]
"00111011110000010000000000100011",	-- 993: 	lw	%r1, [%sp + 35]
"00111100001110110000000000001001",	-- 994: 	sw	%r1, [%r27 + 9]
"00111101001110110000000000001000",	-- 995: 	sw	%r9, [%r27 + 8]
"00111101101110110000000000000111",	-- 996: 	sw	%r13, [%r27 + 7]
"00111011110000010000000000100000",	-- 997: 	lw	%r1, [%sp + 32]
"00111100001110110000000000000110",	-- 998: 	sw	%r1, [%r27 + 6]
"00111101000110110000000000000101",	-- 999: 	sw	%r8, [%r27 + 5]
"00111101010110110000000000000100",	-- 1000: 	sw	%r10, [%r27 + 4]
"00111101111110110000000000000011",	-- 1001: 	sw	%r15, [%r27 + 3]
"00111100110110110000000000000010",	-- 1002: 	sw	%r6, [%r27 + 2]
"00111100010110110000000000000001",	-- 1003: 	sw	%r2, [%r27 + 1]
"11001100000000010000000010000000",	-- 1004: 	lli	%r1, 128
"11001100000000100000000010000000",	-- 1005: 	lli	%r2, 128
"00111111111111100000000000100101",	-- 1006: 	sw	%ra, [%sp + 37]
"00111011011110100000000000000000",	-- 1007: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100110",	-- 1008: 	addi	%sp, %sp, 38
"01010011010000000000000000000000",	-- 1009: 	jalr	%r26
"10101011110111100000000000100110",	-- 1010: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 1011: 	lw	%ra, [%sp + 37]
"11001100000000010000000000000000",	-- 1012: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 1013: 	jr	%ra
	-- halt:
"11111100000000000000000000000000",	-- 1014: 	halt
	-- div10_sub.6209:
"11001100000000110000000000001010",	-- 1015: 	lli	%r3, 10
"00110000011000010000000000000110",	-- 1016: 	bgt	%r3, %r1, bgt_else.8923
"11001100000000110000000000001010",	-- 1017: 	lli	%r3, 10
"10001000001000110000100000000000",	-- 1018: 	sub	%r1, %r1, %r3
"11001100000000110000000000000001",	-- 1019: 	lli	%r3, 1
"10000100010000110001000000000000",	-- 1020: 	add	%r2, %r2, %r3
"01010100000000000000001111110111",	-- 1021: 	j	div10_sub.6209
	-- bgt_else.8923:
"10000100000000100000100000000000",	-- 1022: 	add	%r1, %r0, %r2
"01001111111000000000000000000000",	-- 1023: 	jr	%ra
	-- div10.6193:
"11001100000000100000000000000000",	-- 1024: 	lli	%r2, 0
"01010100000000000000001111110111",	-- 1025: 	j	div10_sub.6209
	-- print_int.2514:
"11001100000000100000000000000000",	-- 1026: 	lli	%r2, 0
"00110000010000010000000000011010",	-- 1027: 	bgt	%r2, %r1, bgt_else.8924
"11001100000000100000000000001010",	-- 1028: 	lli	%r2, 10
"00110000010000010000000000010101",	-- 1029: 	bgt	%r2, %r1, bgt_else.8925
"00111100001111100000000000000000",	-- 1030: 	sw	%r1, [%sp + 0]
"00111111111111100000000000000001",	-- 1031: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 1032: 	addi	%sp, %sp, 2
"01011000000000000000010000000000",	-- 1033: 	jal	div10.6193
"10101011110111100000000000000010",	-- 1034: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 1035: 	lw	%ra, [%sp + 1]
"00111100001111100000000000000001",	-- 1036: 	sw	%r1, [%sp + 1]
"00111111111111100000000000000010",	-- 1037: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1038: 	addi	%sp, %sp, 3
"01011000000000000000010000000010",	-- 1039: 	jal	print_int.2514
"10101011110111100000000000000011",	-- 1040: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1041: 	lw	%ra, [%sp + 2]
"11001100000000010000000000001010",	-- 1042: 	lli	%r1, 10
"00111011110000100000000000000001",	-- 1043: 	lw	%r2, [%sp + 1]
"10001100010000010000100000000000",	-- 1044: 	mul	%r1, %r2, %r1
"00111011110000100000000000000000",	-- 1045: 	lw	%r2, [%sp + 0]
"10001000010000010000100000000000",	-- 1046: 	sub	%r1, %r2, %r1
"11001100000000100000000000110000",	-- 1047: 	lli	%r2, 48
"10000100001000100000100000000000",	-- 1048: 	add	%r1, %r1, %r2
"01010100000000000010101000011010",	-- 1049: 	j	yj_print_char
	-- bgt_else.8925:
"11001100000000100000000000110000",	-- 1050: 	lli	%r2, 48
"10000100001000100000100000000000",	-- 1051: 	add	%r1, %r1, %r2
"01010100000000000010101000011010",	-- 1052: 	j	yj_print_char
	-- bgt_else.8924:
"11001100000000100000000000101101",	-- 1053: 	lli	%r2, 45
"00111100001111100000000000000000",	-- 1054: 	sw	%r1, [%sp + 0]
"10000100000000100000100000000000",	-- 1055: 	add	%r1, %r0, %r2
"00111111111111100000000000000010",	-- 1056: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1057: 	addi	%sp, %sp, 3
"01011000000000000010101000011010",	-- 1058: 	jal	yj_print_char
"10101011110111100000000000000011",	-- 1059: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1060: 	lw	%ra, [%sp + 2]
"00111011110000010000000000000000",	-- 1061: 	lw	%r1, [%sp + 0]
"10001000000000010000100000000000",	-- 1062: 	sub	%r1, %r0, %r1
"01010100000000000000010000000010",	-- 1063: 	j	print_int.2514
	-- calc_sin.6160:
"00010100000000011010101011000001",	-- 1064: 	llif	%f1, -0.166667
"00010000000000011011111000101010",	-- 1065: 	lhif	%f1, -0.166667
"00010100000000101000011100100011",	-- 1066: 	llif	%f2, 0.008333
"00010000000000100011110000001000",	-- 1067: 	lhif	%f2, 0.008333
"00010100000000111001111000111000",	-- 1068: 	llif	%f3, -0.000198
"00010000000000111011100101001111",	-- 1069: 	lhif	%f3, -0.000198
"00010100000001000101001110011100",	-- 1070: 	llif	%f4, 0.000003
"00010000000001000011011001001001",	-- 1071: 	lhif	%f4, 0.000003
"00010100000001010000000000000000",	-- 1072: 	llif	%f5, 0.000000
"00010000000001010000000000000000",	-- 1073: 	lhif	%f5, 0.000000
"00010100000001100000000000000000",	-- 1074: 	llif	%f6, 0.000000
"00010000000001100000000000000000",	-- 1075: 	lhif	%f6, 0.000000
"11101000000000000011100000000000",	-- 1076: 	mulf	%f7, %f0, %f0
"11101000111000000100000000000000",	-- 1077: 	mulf	%f8, %f7, %f0
"11101000111001100011000000000000",	-- 1078: 	mulf	%f6, %f7, %f6
"11100000101001100010100000000000",	-- 1079: 	addf	%f5, %f5, %f6
"11101000111001010010100000000000",	-- 1080: 	mulf	%f5, %f7, %f5
"11100000100001010010000000000000",	-- 1081: 	addf	%f4, %f4, %f5
"11101000111001000010000000000000",	-- 1082: 	mulf	%f4, %f7, %f4
"11100000011001000001100000000000",	-- 1083: 	addf	%f3, %f3, %f4
"11101000111000110001100000000000",	-- 1084: 	mulf	%f3, %f7, %f3
"11100000010000110001000000000000",	-- 1085: 	addf	%f2, %f2, %f3
"11101000111000100001000000000000",	-- 1086: 	mulf	%f2, %f7, %f2
"11100000001000100000100000000000",	-- 1087: 	addf	%f1, %f1, %f2
"11101001000000010000100000000000",	-- 1088: 	mulf	%f1, %f8, %f1
"11100000000000010000000000000000",	-- 1089: 	addf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 1090: 	jr	%ra
	-- sinf__.6162:
"00010100000000010000111111011000",	-- 1091: 	llif	%f1, 1.570796
"00010000000000010011111111001001",	-- 1092: 	lhif	%f1, 1.570796
"00010100000000100000111111011100",	-- 1093: 	llif	%f2, 3.141593
"00010000000000100100000001001001",	-- 1094: 	lhif	%f2, 3.141593
"00010100000000110000111111011010",	-- 1095: 	llif	%f3, 6.283185
"00010000000000110100000011001001",	-- 1096: 	lhif	%f3, 6.283185
"00100000000000110000000000001110",	-- 1097: 	bgtf	%f0, %f3, bgtf_else.8926
"00100000000000100000000000000101",	-- 1098: 	bgtf	%f0, %f2, bgtf_else.8927
"00100000000000010000000000000010",	-- 1099: 	bgtf	%f0, %f1, bgtf_else.8928
"01010100000000000000010000101000",	-- 1100: 	j	calc_sin.6160
	-- bgtf_else.8928:
"11100100010000000000000000000000",	-- 1101: 	subf	%f0, %f2, %f0
"01010100000000000000010001000011",	-- 1102: 	j	sinf__.6162
	-- bgtf_else.8927:
"11100100000000100000000000000000",	-- 1103: 	subf	%f0, %f0, %f2
"00111111111111100000000000000000",	-- 1104: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 1105: 	addi	%sp, %sp, 1
"01011000000000000000010001000011",	-- 1106: 	jal	sinf__.6162
"10101011110111100000000000000001",	-- 1107: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 1108: 	lw	%ra, [%sp + 0]
"00011000000000000000000000000000",	-- 1109: 	negf	%f0, %f0
"01001111111000000000000000000000",	-- 1110: 	jr	%ra
	-- bgtf_else.8926:
"11100100000000110000000000000000",	-- 1111: 	subf	%f0, %f0, %f3
"01010100000000000000010001000011",	-- 1112: 	j	sinf__.6162
	-- sin.2516:
"00010100000000010000000000000000",	-- 1113: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 1114: 	lhif	%f1, 0.000000
"00100000001000000000000000000010",	-- 1115: 	bgtf	%f1, %f0, bgtf_else.8929
"01010100000000000000010001000011",	-- 1116: 	j	sinf__.6162
	-- bgtf_else.8929:
"00011000000000000000000000000000",	-- 1117: 	negf	%f0, %f0
"00111111111111100000000000000000",	-- 1118: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 1119: 	addi	%sp, %sp, 1
"01011000000000000000010001000011",	-- 1120: 	jal	sinf__.6162
"10101011110111100000000000000001",	-- 1121: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 1122: 	lw	%ra, [%sp + 0]
"00011000000000000000000000000000",	-- 1123: 	negf	%f0, %f0
"01001111111000000000000000000000",	-- 1124: 	jr	%ra
	-- calc_cos.6127:
"00010100000000011010101100000100",	-- 1125: 	llif	%f1, 0.041667
"00010000000000010011110100101010",	-- 1126: 	lhif	%f1, 0.041667
"00010100000000100000111100011011",	-- 1127: 	llif	%f2, -0.001389
"00010000000000101011101010110110",	-- 1128: 	lhif	%f2, -0.001389
"00010100000000111011011100010111",	-- 1129: 	llif	%f3, 0.000025
"00010000000000110011011111010001",	-- 1130: 	lhif	%f3, 0.000025
"00010100000001000000000000000000",	-- 1131: 	llif	%f4, -0.000000
"00010000000001001000000000000000",	-- 1132: 	lhif	%f4, -0.000000
"00010100000001010000000000000000",	-- 1133: 	llif	%f5, -0.000000
"00010000000001011000000000000000",	-- 1134: 	lhif	%f5, -0.000000
"11101000000000000000000000000000",	-- 1135: 	mulf	%f0, %f0, %f0
"11101000000001010010100000000000",	-- 1136: 	mulf	%f5, %f0, %f5
"11100000100001010010000000000000",	-- 1137: 	addf	%f4, %f4, %f5
"11101000000001000010000000000000",	-- 1138: 	mulf	%f4, %f0, %f4
"11100000011001000001100000000000",	-- 1139: 	addf	%f3, %f3, %f4
"11101000000000110001100000000000",	-- 1140: 	mulf	%f3, %f0, %f3
"11100000010000110001000000000000",	-- 1141: 	addf	%f2, %f2, %f3
"11101000000000100001000000000000",	-- 1142: 	mulf	%f2, %f0, %f2
"11100000001000100000100000000000",	-- 1143: 	addf	%f1, %f1, %f2
"11101000000000010000100000000000",	-- 1144: 	mulf	%f1, %f0, %f1
"00010100000000100000000000000000",	-- 1145: 	llif	%f2, 1.000000
"00010000000000100011111110000000",	-- 1146: 	lhif	%f2, 1.000000
"00010100000000110000000000000000",	-- 1147: 	llif	%f3, 0.500000
"00010000000000110011111100000000",	-- 1148: 	lhif	%f3, 0.500000
"11101000011000000001100000000000",	-- 1149: 	mulf	%f3, %f3, %f0
"11100100010000110001000000000000",	-- 1150: 	subf	%f2, %f2, %f3
"11101000000000010000000000000000",	-- 1151: 	mulf	%f0, %f0, %f1
"11100000010000000000000000000000",	-- 1152: 	addf	%f0, %f2, %f0
"01001111111000000000000000000000",	-- 1153: 	jr	%ra
	-- cosf__.6129:
"00010100000000010000111111011000",	-- 1154: 	llif	%f1, 1.570796
"00010000000000010011111111001001",	-- 1155: 	lhif	%f1, 1.570796
"00010100000000100000111111011100",	-- 1156: 	llif	%f2, 3.141593
"00010000000000100100000001001001",	-- 1157: 	lhif	%f2, 3.141593
"00010100000000110000111111011010",	-- 1158: 	llif	%f3, 6.283185
"00010000000000110100000011001001",	-- 1159: 	lhif	%f3, 6.283185
"00100000000000110000000000001110",	-- 1160: 	bgtf	%f0, %f3, bgtf_else.8930
"00100000000000100000000000000101",	-- 1161: 	bgtf	%f0, %f2, bgtf_else.8931
"00100000000000010000000000000010",	-- 1162: 	bgtf	%f0, %f1, bgtf_else.8932
"01010100000000000000010001100101",	-- 1163: 	j	calc_cos.6127
	-- bgtf_else.8932:
"11100100010000000000000000000000",	-- 1164: 	subf	%f0, %f2, %f0
"01010100000000000000010010000010",	-- 1165: 	j	cosf__.6129
	-- bgtf_else.8931:
"11100100000000100000000000000000",	-- 1166: 	subf	%f0, %f0, %f2
"00111111111111100000000000000000",	-- 1167: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 1168: 	addi	%sp, %sp, 1
"01011000000000000000010010000010",	-- 1169: 	jal	cosf__.6129
"10101011110111100000000000000001",	-- 1170: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 1171: 	lw	%ra, [%sp + 0]
"00011000000000000000000000000000",	-- 1172: 	negf	%f0, %f0
"01001111111000000000000000000000",	-- 1173: 	jr	%ra
	-- bgtf_else.8930:
"11100100000000110000000000000000",	-- 1174: 	subf	%f0, %f0, %f3
"01010100000000000000010010000010",	-- 1175: 	j	cosf__.6129
	-- cos.2518:
"00010100000000010000000000000000",	-- 1176: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 1177: 	lhif	%f1, 0.000000
"00100000001000000000000000000010",	-- 1178: 	bgtf	%f1, %f0, bgtf_else.8933
"01010100000000000000010010000010",	-- 1179: 	j	cosf__.6129
	-- bgtf_else.8933:
"00011000000000000000000000000000",	-- 1180: 	negf	%f0, %f0
"01010100000000000000010010000010",	-- 1181: 	j	cosf__.6129
	-- atan.2520:
"10110000000111100000000000000000",	-- 1182: 	sf	%f0, [%sp + 0]
"00111111111111100000000000000001",	-- 1183: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 1184: 	addi	%sp, %sp, 2
"01011000000000000010101001001111",	-- 1185: 	jal	yj_fabs
"10101011110111100000000000000010",	-- 1186: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 1187: 	lw	%ra, [%sp + 1]
"00010100000000011001100110011010",	-- 1188: 	llif	%f1, 0.150000
"00010000000000010011111000011001",	-- 1189: 	lhif	%f1, 0.150000
"00100000000000010000000000010011",	-- 1190: 	bgtf	%f0, %f1, bgtf_else.8934
"10010011110000000000000000000000",	-- 1191: 	lf	%f0, [%sp + 0]
"11101000000000000000100000000000",	-- 1192: 	mulf	%f1, %f0, %f0
"00010100000000100000000000000000",	-- 1193: 	llif	%f2, 1.000000
"00010000000000100011111110000000",	-- 1194: 	lhif	%f2, 1.000000
"00010100000000111010101010011111",	-- 1195: 	llif	%f3, -0.333333
"00010000000000111011111010101010",	-- 1196: 	lhif	%f3, -0.333333
"00010100000001001100110011001101",	-- 1197: 	llif	%f4, 0.200000
"00010000000001000011111001001100",	-- 1198: 	lhif	%f4, 0.200000
"00010100000001010100100100011011",	-- 1199: 	llif	%f5, 0.142857
"00010000000001010011111000010010",	-- 1200: 	lhif	%f5, 0.142857
"11101000001001010010100000000000",	-- 1201: 	mulf	%f5, %f1, %f5
"11100000100001010010000000000000",	-- 1202: 	addf	%f4, %f4, %f5
"11101000001001000010000000000000",	-- 1203: 	mulf	%f4, %f1, %f4
"11100000011001000001100000000000",	-- 1204: 	addf	%f3, %f3, %f4
"11101000001000110000100000000000",	-- 1205: 	mulf	%f1, %f1, %f3
"11100000010000010000100000000000",	-- 1206: 	addf	%f1, %f2, %f1
"11101000000000010000000000000000",	-- 1207: 	mulf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 1208: 	jr	%ra
	-- bgtf_else.8934:
"00010100000000000000000000000000",	-- 1209: 	llif	%f0, -1.000000
"00010000000000001011111110000000",	-- 1210: 	lhif	%f0, -1.000000
"00010100000000010000000000000000",	-- 1211: 	llif	%f1, 1.000000
"00010000000000010011111110000000",	-- 1212: 	lhif	%f1, 1.000000
"10010011110000100000000000000000",	-- 1213: 	lf	%f2, [%sp + 0]
"11101000010000100001100000000000",	-- 1214: 	mulf	%f3, %f2, %f2
"11100000001000110000100000000000",	-- 1215: 	addf	%f1, %f1, %f3
"10110000000111100000000000000001",	-- 1216: 	sf	%f0, [%sp + 1]
"00001100001000000000000000000000",	-- 1217: 	movf	%f0, %f1
"00111111111111100000000000000010",	-- 1218: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1219: 	addi	%sp, %sp, 3
"01011000000000000010101000110000",	-- 1220: 	jal	yj_sqrt
"10101011110111100000000000000011",	-- 1221: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1222: 	lw	%ra, [%sp + 2]
"10010011110000010000000000000001",	-- 1223: 	lf	%f1, [%sp + 1]
"11100000001000000000000000000000",	-- 1224: 	addf	%f0, %f1, %f0
"10010011110000010000000000000000",	-- 1225: 	lf	%f1, [%sp + 0]
"11101100000000010000000000000000",	-- 1226: 	divf	%f0, %f0, %f1
"00010100000000010000000000000000",	-- 1227: 	llif	%f1, 2.000000
"00010000000000010100000000000000",	-- 1228: 	lhif	%f1, 2.000000
"10110000001111100000000000000010",	-- 1229: 	sf	%f1, [%sp + 2]
"00111111111111100000000000000011",	-- 1230: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 1231: 	addi	%sp, %sp, 4
"01011000000000000000010010011110",	-- 1232: 	jal	atan.2520
"10101011110111100000000000000100",	-- 1233: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 1234: 	lw	%ra, [%sp + 3]
"10010011110000010000000000000010",	-- 1235: 	lf	%f1, [%sp + 2]
"11101000001000000000000000000000",	-- 1236: 	mulf	%f0, %f1, %f0
"01001111111000000000000000000000",	-- 1237: 	jr	%ra
	-- fispos.2522:
"00010100000000010000000000000000",	-- 1238: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 1239: 	lhif	%f1, 0.000000
"00100000000000010000000000000011",	-- 1240: 	bgtf	%f0, %f1, bgtf_else.8935
"11001100000000010000000000000000",	-- 1241: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 1242: 	jr	%ra
	-- bgtf_else.8935:
"11001100000000010000000000000001",	-- 1243: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 1244: 	jr	%ra
	-- fisneg.2524:
"00010100000000010000000000000000",	-- 1245: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 1246: 	lhif	%f1, 0.000000
"00100000001000000000000000000011",	-- 1247: 	bgtf	%f1, %f0, bgtf_else.8936
"11001100000000010000000000000000",	-- 1248: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 1249: 	jr	%ra
	-- bgtf_else.8936:
"11001100000000010000000000000001",	-- 1250: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 1251: 	jr	%ra
	-- fiszero.2526:
"00010100000000010000000000000000",	-- 1252: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 1253: 	lhif	%f1, 0.000000
"01011100000000010000000000000000",	-- 1254: 	movf2i	%r1, %f0
"01011100001000100000000000000000",	-- 1255: 	movf2i	%r2, %f1
"00101000001000100000000000000011",	-- 1256: 	bneq	%r1, %r2, bneq_else.8937
"11001100000000010000000000000001",	-- 1257: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 1258: 	jr	%ra
	-- bneq_else.8937:
"11001100000000010000000000000000",	-- 1259: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 1260: 	jr	%ra
	-- fhalf.2528:
"00010100000000010000000000000000",	-- 1261: 	llif	%f1, 0.500000
"00010000000000010011111100000000",	-- 1262: 	lhif	%f1, 0.500000
"11101000000000010000000000000000",	-- 1263: 	mulf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 1264: 	jr	%ra
	-- fsqr.2530:
"11101000000000000000000000000000",	-- 1265: 	mulf	%f0, %f0, %f0
"01001111111000000000000000000000",	-- 1266: 	jr	%ra
	-- fless.2532:
"00100000001000000000000000000011",	-- 1267: 	bgtf	%f1, %f0, bgtf_else.8938
"11001100000000010000000000000000",	-- 1268: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 1269: 	jr	%ra
	-- bgtf_else.8938:
"11001100000000010000000000000001",	-- 1270: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 1271: 	jr	%ra
	-- xor.2565:
"11001100000000110000000000000000",	-- 1272: 	lli	%r3, 0
"00101000001000110000000000000011",	-- 1273: 	bneq	%r1, %r3, bneq_else.8939
"10000100000000100000100000000000",	-- 1274: 	add	%r1, %r0, %r2
"01001111111000000000000000000000",	-- 1275: 	jr	%ra
	-- bneq_else.8939:
"11001100000000010000000000000000",	-- 1276: 	lli	%r1, 0
"00101000010000010000000000000011",	-- 1277: 	bneq	%r2, %r1, bneq_else.8940
"11001100000000010000000000000001",	-- 1278: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 1279: 	jr	%ra
	-- bneq_else.8940:
"11001100000000010000000000000000",	-- 1280: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 1281: 	jr	%ra
	-- sgn.2568:
"10110000000111100000000000000000",	-- 1282: 	sf	%f0, [%sp + 0]
"00111111111111100000000000000001",	-- 1283: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 1284: 	addi	%sp, %sp, 2
"01011000000000000000010011100100",	-- 1285: 	jal	fiszero.2526
"10101011110111100000000000000010",	-- 1286: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 1287: 	lw	%ra, [%sp + 1]
"11001100000000100000000000000000",	-- 1288: 	lli	%r2, 0
"00101000001000100000000000001111",	-- 1289: 	bneq	%r1, %r2, bneq_else.8941
"10010011110000000000000000000000",	-- 1290: 	lf	%f0, [%sp + 0]
"00111111111111100000000000000001",	-- 1291: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 1292: 	addi	%sp, %sp, 2
"01011000000000000000010011010110",	-- 1293: 	jal	fispos.2522
"10101011110111100000000000000010",	-- 1294: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 1295: 	lw	%ra, [%sp + 1]
"11001100000000100000000000000000",	-- 1296: 	lli	%r2, 0
"00101000001000100000000000000100",	-- 1297: 	bneq	%r1, %r2, bneq_else.8942
"00010100000000000000000000000000",	-- 1298: 	llif	%f0, -1.000000
"00010000000000001011111110000000",	-- 1299: 	lhif	%f0, -1.000000
"01001111111000000000000000000000",	-- 1300: 	jr	%ra
	-- bneq_else.8942:
"00010100000000000000000000000000",	-- 1301: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 1302: 	lhif	%f0, 1.000000
"01001111111000000000000000000000",	-- 1303: 	jr	%ra
	-- bneq_else.8941:
"00010100000000000000000000000000",	-- 1304: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 1305: 	lhif	%f0, 0.000000
"01001111111000000000000000000000",	-- 1306: 	jr	%ra
	-- fneg_cond.2570:
"11001100000000100000000000000000",	-- 1307: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 1308: 	bneq	%r1, %r2, bneq_else.8943
"01010100000000000010101001010001",	-- 1309: 	j	yj_fneg
	-- bneq_else.8943:
"01001111111000000000000000000000",	-- 1310: 	jr	%ra
	-- add_mod5.2573:
"10000100001000100000100000000000",	-- 1311: 	add	%r1, %r1, %r2
"11001100000000100000000000000101",	-- 1312: 	lli	%r2, 5
"00110000010000010000000000000100",	-- 1313: 	bgt	%r2, %r1, bgt_else.8944
"11001100000000100000000000000101",	-- 1314: 	lli	%r2, 5
"10001000001000100000100000000000",	-- 1315: 	sub	%r1, %r1, %r2
"01001111111000000000000000000000",	-- 1316: 	jr	%ra
	-- bgt_else.8944:
"01001111111000000000000000000000",	-- 1317: 	jr	%ra
	-- vecset.2576:
"11001100000000100000000000000000",	-- 1318: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 1319: 	add	%r2, %r1, %r2
"10110000000000100000000000000000",	-- 1320: 	sf	%f0, [%r2 + 0]
"11001100000000100000000000000001",	-- 1321: 	lli	%r2, 1
"10000100001000100001000000000000",	-- 1322: 	add	%r2, %r1, %r2
"10110000001000100000000000000000",	-- 1323: 	sf	%f1, [%r2 + 0]
"11001100000000100000000000000010",	-- 1324: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1325: 	add	%r1, %r1, %r2
"10110000010000010000000000000000",	-- 1326: 	sf	%f2, [%r1 + 0]
"01001111111000000000000000000000",	-- 1327: 	jr	%ra
	-- vecfill.2581:
"11001100000000100000000000000000",	-- 1328: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 1329: 	add	%r2, %r1, %r2
"10110000000000100000000000000000",	-- 1330: 	sf	%f0, [%r2 + 0]
"11001100000000100000000000000001",	-- 1331: 	lli	%r2, 1
"10000100001000100001000000000000",	-- 1332: 	add	%r2, %r1, %r2
"10110000000000100000000000000000",	-- 1333: 	sf	%f0, [%r2 + 0]
"11001100000000100000000000000010",	-- 1334: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1335: 	add	%r1, %r1, %r2
"10110000000000010000000000000000",	-- 1336: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1337: 	jr	%ra
	-- vecbzero.2584:
"00010100000000000000000000000000",	-- 1338: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 1339: 	lhif	%f0, 0.000000
"01010100000000000000010100110000",	-- 1340: 	j	vecfill.2581
	-- veccpy.2586:
"11001100000000110000000000000000",	-- 1341: 	lli	%r3, 0
"11001100000001000000000000000000",	-- 1342: 	lli	%r4, 0
"10000100010001000010000000000000",	-- 1343: 	add	%r4, %r2, %r4
"10010000100000000000000000000000",	-- 1344: 	lf	%f0, [%r4 + 0]
"10000100001000110001100000000000",	-- 1345: 	add	%r3, %r1, %r3
"10110000000000110000000000000000",	-- 1346: 	sf	%f0, [%r3 + 0]
"11001100000000110000000000000001",	-- 1347: 	lli	%r3, 1
"11001100000001000000000000000001",	-- 1348: 	lli	%r4, 1
"10000100010001000010000000000000",	-- 1349: 	add	%r4, %r2, %r4
"10010000100000000000000000000000",	-- 1350: 	lf	%f0, [%r4 + 0]
"10000100001000110001100000000000",	-- 1351: 	add	%r3, %r1, %r3
"10110000000000110000000000000000",	-- 1352: 	sf	%f0, [%r3 + 0]
"11001100000000110000000000000010",	-- 1353: 	lli	%r3, 2
"11001100000001000000000000000010",	-- 1354: 	lli	%r4, 2
"10000100010001000001000000000000",	-- 1355: 	add	%r2, %r2, %r4
"10010000010000000000000000000000",	-- 1356: 	lf	%f0, [%r2 + 0]
"10000100001000110000100000000000",	-- 1357: 	add	%r1, %r1, %r3
"10110000000000010000000000000000",	-- 1358: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1359: 	jr	%ra
	-- vecunit_sgn.2594:
"11001100000000110000000000000000",	-- 1360: 	lli	%r3, 0
"10000100001000110001100000000000",	-- 1361: 	add	%r3, %r1, %r3
"10010000011000000000000000000000",	-- 1362: 	lf	%f0, [%r3 + 0]
"00111100010111100000000000000000",	-- 1363: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 1364: 	sw	%r1, [%sp + 1]
"00111111111111100000000000000010",	-- 1365: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1366: 	addi	%sp, %sp, 3
"01011000000000000000010011110001",	-- 1367: 	jal	fsqr.2530
"10101011110111100000000000000011",	-- 1368: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1369: 	lw	%ra, [%sp + 2]
"11001100000000010000000000000001",	-- 1370: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 1371: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 1372: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 1373: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000010",	-- 1374: 	sf	%f0, [%sp + 2]
"00001100001000000000000000000000",	-- 1375: 	movf	%f0, %f1
"00111111111111100000000000000011",	-- 1376: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 1377: 	addi	%sp, %sp, 4
"01011000000000000000010011110001",	-- 1378: 	jal	fsqr.2530
"10101011110111100000000000000100",	-- 1379: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 1380: 	lw	%ra, [%sp + 3]
"10010011110000010000000000000010",	-- 1381: 	lf	%f1, [%sp + 2]
"11100000001000000000000000000000",	-- 1382: 	addf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 1383: 	lli	%r1, 2
"00111011110000100000000000000001",	-- 1384: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 1385: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 1386: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000011",	-- 1387: 	sf	%f0, [%sp + 3]
"00001100001000000000000000000000",	-- 1388: 	movf	%f0, %f1
"00111111111111100000000000000100",	-- 1389: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 1390: 	addi	%sp, %sp, 5
"01011000000000000000010011110001",	-- 1391: 	jal	fsqr.2530
"10101011110111100000000000000101",	-- 1392: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 1393: 	lw	%ra, [%sp + 4]
"10010011110000010000000000000011",	-- 1394: 	lf	%f1, [%sp + 3]
"11100000001000000000000000000000",	-- 1395: 	addf	%f0, %f1, %f0
"00111111111111100000000000000100",	-- 1396: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 1397: 	addi	%sp, %sp, 5
"01011000000000000010101000110000",	-- 1398: 	jal	yj_sqrt
"10101011110111100000000000000101",	-- 1399: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 1400: 	lw	%ra, [%sp + 4]
"10110000000111100000000000000100",	-- 1401: 	sf	%f0, [%sp + 4]
"00111111111111100000000000000101",	-- 1402: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 1403: 	addi	%sp, %sp, 6
"01011000000000000000010011100100",	-- 1404: 	jal	fiszero.2526
"10101011110111100000000000000110",	-- 1405: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 1406: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000000",	-- 1407: 	lli	%r2, 0
"00101000001000100000000000001110",	-- 1408: 	bneq	%r1, %r2, bneq_else.8948
"11001100000000010000000000000000",	-- 1409: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 1410: 	lw	%r2, [%sp + 0]
"00101000010000010000000000000110",	-- 1411: 	bneq	%r2, %r1, bneq_else.8950
"00010100000000000000000000000000",	-- 1412: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 1413: 	lhif	%f0, 1.000000
"10010011110000010000000000000100",	-- 1414: 	lf	%f1, [%sp + 4]
"11101100000000010000000000000000",	-- 1415: 	divf	%f0, %f0, %f1
"01010100000000000000010110001101",	-- 1416: 	j	bneq_cont.8951
	-- bneq_else.8950:
"00010100000000000000000000000000",	-- 1417: 	llif	%f0, -1.000000
"00010000000000001011111110000000",	-- 1418: 	lhif	%f0, -1.000000
"10010011110000010000000000000100",	-- 1419: 	lf	%f1, [%sp + 4]
"11101100000000010000000000000000",	-- 1420: 	divf	%f0, %f0, %f1
	-- bneq_cont.8951:
"01010100000000000000010110010000",	-- 1421: 	j	bneq_cont.8949
	-- bneq_else.8948:
"00010100000000000000000000000000",	-- 1422: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 1423: 	lhif	%f0, 1.000000
	-- bneq_cont.8949:
"11001100000000010000000000000000",	-- 1424: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 1425: 	lli	%r2, 0
"00111011110000110000000000000001",	-- 1426: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 1427: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 1428: 	lf	%f1, [%r2 + 0]
"11101000001000000000100000000000",	-- 1429: 	mulf	%f1, %f1, %f0
"10000100011000010000100000000000",	-- 1430: 	add	%r1, %r3, %r1
"10110000001000010000000000000000",	-- 1431: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000001",	-- 1432: 	lli	%r1, 1
"11001100000000100000000000000001",	-- 1433: 	lli	%r2, 1
"10000100011000100001000000000000",	-- 1434: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 1435: 	lf	%f1, [%r2 + 0]
"11101000001000000000100000000000",	-- 1436: 	mulf	%f1, %f1, %f0
"10000100011000010000100000000000",	-- 1437: 	add	%r1, %r3, %r1
"10110000001000010000000000000000",	-- 1438: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 1439: 	lli	%r1, 2
"11001100000000100000000000000010",	-- 1440: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 1441: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 1442: 	lf	%f1, [%r2 + 0]
"11101000001000000000000000000000",	-- 1443: 	mulf	%f0, %f1, %f0
"10000100011000010000100000000000",	-- 1444: 	add	%r1, %r3, %r1
"10110000000000010000000000000000",	-- 1445: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1446: 	jr	%ra
	-- veciprod.2597:
"11001100000000110000000000000000",	-- 1447: 	lli	%r3, 0
"10000100001000110001100000000000",	-- 1448: 	add	%r3, %r1, %r3
"10010000011000000000000000000000",	-- 1449: 	lf	%f0, [%r3 + 0]
"11001100000000110000000000000000",	-- 1450: 	lli	%r3, 0
"10000100010000110001100000000000",	-- 1451: 	add	%r3, %r2, %r3
"10010000011000010000000000000000",	-- 1452: 	lf	%f1, [%r3 + 0]
"11101000000000010000000000000000",	-- 1453: 	mulf	%f0, %f0, %f1
"11001100000000110000000000000001",	-- 1454: 	lli	%r3, 1
"10000100001000110001100000000000",	-- 1455: 	add	%r3, %r1, %r3
"10010000011000010000000000000000",	-- 1456: 	lf	%f1, [%r3 + 0]
"11001100000000110000000000000001",	-- 1457: 	lli	%r3, 1
"10000100010000110001100000000000",	-- 1458: 	add	%r3, %r2, %r3
"10010000011000100000000000000000",	-- 1459: 	lf	%f2, [%r3 + 0]
"11101000001000100000100000000000",	-- 1460: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 1461: 	addf	%f0, %f0, %f1
"11001100000000110000000000000010",	-- 1462: 	lli	%r3, 2
"10000100001000110000100000000000",	-- 1463: 	add	%r1, %r1, %r3
"10010000001000010000000000000000",	-- 1464: 	lf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 1465: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 1466: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 1467: 	lf	%f2, [%r1 + 0]
"11101000001000100000100000000000",	-- 1468: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 1469: 	addf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 1470: 	jr	%ra
	-- veciprod2.2600:
"11001100000000100000000000000000",	-- 1471: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 1472: 	add	%r2, %r1, %r2
"10010000010000110000000000000000",	-- 1473: 	lf	%f3, [%r2 + 0]
"11101000011000000000000000000000",	-- 1474: 	mulf	%f0, %f3, %f0
"11001100000000100000000000000001",	-- 1475: 	lli	%r2, 1
"10000100001000100001000000000000",	-- 1476: 	add	%r2, %r1, %r2
"10010000010000110000000000000000",	-- 1477: 	lf	%f3, [%r2 + 0]
"11101000011000010000100000000000",	-- 1478: 	mulf	%f1, %f3, %f1
"11100000000000010000000000000000",	-- 1479: 	addf	%f0, %f0, %f1
"11001100000000100000000000000010",	-- 1480: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1481: 	add	%r1, %r1, %r2
"10010000001000010000000000000000",	-- 1482: 	lf	%f1, [%r1 + 0]
"11101000001000100000100000000000",	-- 1483: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 1484: 	addf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 1485: 	jr	%ra
	-- vecaccum.2605:
"11001100000000110000000000000000",	-- 1486: 	lli	%r3, 0
"11001100000001000000000000000000",	-- 1487: 	lli	%r4, 0
"10000100001001000010000000000000",	-- 1488: 	add	%r4, %r1, %r4
"10010000100000010000000000000000",	-- 1489: 	lf	%f1, [%r4 + 0]
"11001100000001000000000000000000",	-- 1490: 	lli	%r4, 0
"10000100010001000010000000000000",	-- 1491: 	add	%r4, %r2, %r4
"10010000100000100000000000000000",	-- 1492: 	lf	%f2, [%r4 + 0]
"11101000000000100001000000000000",	-- 1493: 	mulf	%f2, %f0, %f2
"11100000001000100000100000000000",	-- 1494: 	addf	%f1, %f1, %f2
"10000100001000110001100000000000",	-- 1495: 	add	%r3, %r1, %r3
"10110000001000110000000000000000",	-- 1496: 	sf	%f1, [%r3 + 0]
"11001100000000110000000000000001",	-- 1497: 	lli	%r3, 1
"11001100000001000000000000000001",	-- 1498: 	lli	%r4, 1
"10000100001001000010000000000000",	-- 1499: 	add	%r4, %r1, %r4
"10010000100000010000000000000000",	-- 1500: 	lf	%f1, [%r4 + 0]
"11001100000001000000000000000001",	-- 1501: 	lli	%r4, 1
"10000100010001000010000000000000",	-- 1502: 	add	%r4, %r2, %r4
"10010000100000100000000000000000",	-- 1503: 	lf	%f2, [%r4 + 0]
"11101000000000100001000000000000",	-- 1504: 	mulf	%f2, %f0, %f2
"11100000001000100000100000000000",	-- 1505: 	addf	%f1, %f1, %f2
"10000100001000110001100000000000",	-- 1506: 	add	%r3, %r1, %r3
"10110000001000110000000000000000",	-- 1507: 	sf	%f1, [%r3 + 0]
"11001100000000110000000000000010",	-- 1508: 	lli	%r3, 2
"11001100000001000000000000000010",	-- 1509: 	lli	%r4, 2
"10000100001001000010000000000000",	-- 1510: 	add	%r4, %r1, %r4
"10010000100000010000000000000000",	-- 1511: 	lf	%f1, [%r4 + 0]
"11001100000001000000000000000010",	-- 1512: 	lli	%r4, 2
"10000100010001000001000000000000",	-- 1513: 	add	%r2, %r2, %r4
"10010000010000100000000000000000",	-- 1514: 	lf	%f2, [%r2 + 0]
"11101000000000100000000000000000",	-- 1515: 	mulf	%f0, %f0, %f2
"11100000001000000000000000000000",	-- 1516: 	addf	%f0, %f1, %f0
"10000100001000110000100000000000",	-- 1517: 	add	%r1, %r1, %r3
"10110000000000010000000000000000",	-- 1518: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1519: 	jr	%ra
	-- vecadd.2609:
"11001100000000110000000000000000",	-- 1520: 	lli	%r3, 0
"11001100000001000000000000000000",	-- 1521: 	lli	%r4, 0
"10000100001001000010000000000000",	-- 1522: 	add	%r4, %r1, %r4
"10010000100000000000000000000000",	-- 1523: 	lf	%f0, [%r4 + 0]
"11001100000001000000000000000000",	-- 1524: 	lli	%r4, 0
"10000100010001000010000000000000",	-- 1525: 	add	%r4, %r2, %r4
"10010000100000010000000000000000",	-- 1526: 	lf	%f1, [%r4 + 0]
"11100000000000010000000000000000",	-- 1527: 	addf	%f0, %f0, %f1
"10000100001000110001100000000000",	-- 1528: 	add	%r3, %r1, %r3
"10110000000000110000000000000000",	-- 1529: 	sf	%f0, [%r3 + 0]
"11001100000000110000000000000001",	-- 1530: 	lli	%r3, 1
"11001100000001000000000000000001",	-- 1531: 	lli	%r4, 1
"10000100001001000010000000000000",	-- 1532: 	add	%r4, %r1, %r4
"10010000100000000000000000000000",	-- 1533: 	lf	%f0, [%r4 + 0]
"11001100000001000000000000000001",	-- 1534: 	lli	%r4, 1
"10000100010001000010000000000000",	-- 1535: 	add	%r4, %r2, %r4
"10010000100000010000000000000000",	-- 1536: 	lf	%f1, [%r4 + 0]
"11100000000000010000000000000000",	-- 1537: 	addf	%f0, %f0, %f1
"10000100001000110001100000000000",	-- 1538: 	add	%r3, %r1, %r3
"10110000000000110000000000000000",	-- 1539: 	sf	%f0, [%r3 + 0]
"11001100000000110000000000000010",	-- 1540: 	lli	%r3, 2
"11001100000001000000000000000010",	-- 1541: 	lli	%r4, 2
"10000100001001000010000000000000",	-- 1542: 	add	%r4, %r1, %r4
"10010000100000000000000000000000",	-- 1543: 	lf	%f0, [%r4 + 0]
"11001100000001000000000000000010",	-- 1544: 	lli	%r4, 2
"10000100010001000001000000000000",	-- 1545: 	add	%r2, %r2, %r4
"10010000010000010000000000000000",	-- 1546: 	lf	%f1, [%r2 + 0]
"11100000000000010000000000000000",	-- 1547: 	addf	%f0, %f0, %f1
"10000100001000110000100000000000",	-- 1548: 	add	%r1, %r1, %r3
"10110000000000010000000000000000",	-- 1549: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1550: 	jr	%ra
	-- vecscale.2615:
"11001100000000100000000000000000",	-- 1551: 	lli	%r2, 0
"11001100000000110000000000000000",	-- 1552: 	lli	%r3, 0
"10000100001000110001100000000000",	-- 1553: 	add	%r3, %r1, %r3
"10010000011000010000000000000000",	-- 1554: 	lf	%f1, [%r3 + 0]
"11101000001000000000100000000000",	-- 1555: 	mulf	%f1, %f1, %f0
"10000100001000100001000000000000",	-- 1556: 	add	%r2, %r1, %r2
"10110000001000100000000000000000",	-- 1557: 	sf	%f1, [%r2 + 0]
"11001100000000100000000000000001",	-- 1558: 	lli	%r2, 1
"11001100000000110000000000000001",	-- 1559: 	lli	%r3, 1
"10000100001000110001100000000000",	-- 1560: 	add	%r3, %r1, %r3
"10010000011000010000000000000000",	-- 1561: 	lf	%f1, [%r3 + 0]
"11101000001000000000100000000000",	-- 1562: 	mulf	%f1, %f1, %f0
"10000100001000100001000000000000",	-- 1563: 	add	%r2, %r1, %r2
"10110000001000100000000000000000",	-- 1564: 	sf	%f1, [%r2 + 0]
"11001100000000100000000000000010",	-- 1565: 	lli	%r2, 2
"11001100000000110000000000000010",	-- 1566: 	lli	%r3, 2
"10000100001000110001100000000000",	-- 1567: 	add	%r3, %r1, %r3
"10010000011000010000000000000000",	-- 1568: 	lf	%f1, [%r3 + 0]
"11101000001000000000000000000000",	-- 1569: 	mulf	%f0, %f1, %f0
"10000100001000100000100000000000",	-- 1570: 	add	%r1, %r1, %r2
"10110000000000010000000000000000",	-- 1571: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1572: 	jr	%ra
	-- vecaccumv.2618:
"11001100000001000000000000000000",	-- 1573: 	lli	%r4, 0
"11001100000001010000000000000000",	-- 1574: 	lli	%r5, 0
"10000100001001010010100000000000",	-- 1575: 	add	%r5, %r1, %r5
"10010000101000000000000000000000",	-- 1576: 	lf	%f0, [%r5 + 0]
"11001100000001010000000000000000",	-- 1577: 	lli	%r5, 0
"10000100010001010010100000000000",	-- 1578: 	add	%r5, %r2, %r5
"10010000101000010000000000000000",	-- 1579: 	lf	%f1, [%r5 + 0]
"11001100000001010000000000000000",	-- 1580: 	lli	%r5, 0
"10000100011001010010100000000000",	-- 1581: 	add	%r5, %r3, %r5
"10010000101000100000000000000000",	-- 1582: 	lf	%f2, [%r5 + 0]
"11101000001000100000100000000000",	-- 1583: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 1584: 	addf	%f0, %f0, %f1
"10000100001001000010000000000000",	-- 1585: 	add	%r4, %r1, %r4
"10110000000001000000000000000000",	-- 1586: 	sf	%f0, [%r4 + 0]
"11001100000001000000000000000001",	-- 1587: 	lli	%r4, 1
"11001100000001010000000000000001",	-- 1588: 	lli	%r5, 1
"10000100001001010010100000000000",	-- 1589: 	add	%r5, %r1, %r5
"10010000101000000000000000000000",	-- 1590: 	lf	%f0, [%r5 + 0]
"11001100000001010000000000000001",	-- 1591: 	lli	%r5, 1
"10000100010001010010100000000000",	-- 1592: 	add	%r5, %r2, %r5
"10010000101000010000000000000000",	-- 1593: 	lf	%f1, [%r5 + 0]
"11001100000001010000000000000001",	-- 1594: 	lli	%r5, 1
"10000100011001010010100000000000",	-- 1595: 	add	%r5, %r3, %r5
"10010000101000100000000000000000",	-- 1596: 	lf	%f2, [%r5 + 0]
"11101000001000100000100000000000",	-- 1597: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 1598: 	addf	%f0, %f0, %f1
"10000100001001000010000000000000",	-- 1599: 	add	%r4, %r1, %r4
"10110000000001000000000000000000",	-- 1600: 	sf	%f0, [%r4 + 0]
"11001100000001000000000000000010",	-- 1601: 	lli	%r4, 2
"11001100000001010000000000000010",	-- 1602: 	lli	%r5, 2
"10000100001001010010100000000000",	-- 1603: 	add	%r5, %r1, %r5
"10010000101000000000000000000000",	-- 1604: 	lf	%f0, [%r5 + 0]
"11001100000001010000000000000010",	-- 1605: 	lli	%r5, 2
"10000100010001010001000000000000",	-- 1606: 	add	%r2, %r2, %r5
"10010000010000010000000000000000",	-- 1607: 	lf	%f1, [%r2 + 0]
"11001100000000100000000000000010",	-- 1608: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 1609: 	add	%r2, %r3, %r2
"10010000010000100000000000000000",	-- 1610: 	lf	%f2, [%r2 + 0]
"11101000001000100000100000000000",	-- 1611: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 1612: 	addf	%f0, %f0, %f1
"10000100001001000000100000000000",	-- 1613: 	add	%r1, %r1, %r4
"10110000000000010000000000000000",	-- 1614: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1615: 	jr	%ra
	-- o_texturetype.2622:
"00111000001000010000000000000000",	-- 1616: 	lw	%r1, [%r1 + 0]
"01001111111000000000000000000000",	-- 1617: 	jr	%ra
	-- o_form.2624:
"00111000001000010000000000000001",	-- 1618: 	lw	%r1, [%r1 + 1]
"01001111111000000000000000000000",	-- 1619: 	jr	%ra
	-- o_reflectiontype.2626:
"00111000001000010000000000000010",	-- 1620: 	lw	%r1, [%r1 + 2]
"01001111111000000000000000000000",	-- 1621: 	jr	%ra
	-- o_isinvert.2628:
"00111000001000010000000000000110",	-- 1622: 	lw	%r1, [%r1 + 6]
"01001111111000000000000000000000",	-- 1623: 	jr	%ra
	-- o_isrot.2630:
"00111000001000010000000000000011",	-- 1624: 	lw	%r1, [%r1 + 3]
"01001111111000000000000000000000",	-- 1625: 	jr	%ra
	-- o_param_a.2632:
"00111000001000010000000000000100",	-- 1626: 	lw	%r1, [%r1 + 4]
"11001100000000100000000000000000",	-- 1627: 	lli	%r2, 0
"10000100001000100000100000000000",	-- 1628: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1629: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1630: 	jr	%ra
	-- o_param_b.2634:
"00111000001000010000000000000100",	-- 1631: 	lw	%r1, [%r1 + 4]
"11001100000000100000000000000001",	-- 1632: 	lli	%r2, 1
"10000100001000100000100000000000",	-- 1633: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1634: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1635: 	jr	%ra
	-- o_param_c.2636:
"00111000001000010000000000000100",	-- 1636: 	lw	%r1, [%r1 + 4]
"11001100000000100000000000000010",	-- 1637: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1638: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1639: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1640: 	jr	%ra
	-- o_param_abc.2638:
"00111000001000010000000000000100",	-- 1641: 	lw	%r1, [%r1 + 4]
"01001111111000000000000000000000",	-- 1642: 	jr	%ra
	-- o_param_x.2640:
"00111000001000010000000000000101",	-- 1643: 	lw	%r1, [%r1 + 5]
"11001100000000100000000000000000",	-- 1644: 	lli	%r2, 0
"10000100001000100000100000000000",	-- 1645: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1646: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1647: 	jr	%ra
	-- o_param_y.2642:
"00111000001000010000000000000101",	-- 1648: 	lw	%r1, [%r1 + 5]
"11001100000000100000000000000001",	-- 1649: 	lli	%r2, 1
"10000100001000100000100000000000",	-- 1650: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1651: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1652: 	jr	%ra
	-- o_param_z.2644:
"00111000001000010000000000000101",	-- 1653: 	lw	%r1, [%r1 + 5]
"11001100000000100000000000000010",	-- 1654: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1655: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1656: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1657: 	jr	%ra
	-- o_diffuse.2646:
"00111000001000010000000000000111",	-- 1658: 	lw	%r1, [%r1 + 7]
"11001100000000100000000000000000",	-- 1659: 	lli	%r2, 0
"10000100001000100000100000000000",	-- 1660: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1661: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1662: 	jr	%ra
	-- o_hilight.2648:
"00111000001000010000000000000111",	-- 1663: 	lw	%r1, [%r1 + 7]
"11001100000000100000000000000001",	-- 1664: 	lli	%r2, 1
"10000100001000100000100000000000",	-- 1665: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1666: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1667: 	jr	%ra
	-- o_color_red.2650:
"00111000001000010000000000001000",	-- 1668: 	lw	%r1, [%r1 + 8]
"11001100000000100000000000000000",	-- 1669: 	lli	%r2, 0
"10000100001000100000100000000000",	-- 1670: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1671: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1672: 	jr	%ra
	-- o_color_green.2652:
"00111000001000010000000000001000",	-- 1673: 	lw	%r1, [%r1 + 8]
"11001100000000100000000000000001",	-- 1674: 	lli	%r2, 1
"10000100001000100000100000000000",	-- 1675: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1676: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1677: 	jr	%ra
	-- o_color_blue.2654:
"00111000001000010000000000001000",	-- 1678: 	lw	%r1, [%r1 + 8]
"11001100000000100000000000000010",	-- 1679: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1680: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1681: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1682: 	jr	%ra
	-- o_param_r1.2656:
"00111000001000010000000000001001",	-- 1683: 	lw	%r1, [%r1 + 9]
"11001100000000100000000000000000",	-- 1684: 	lli	%r2, 0
"10000100001000100000100000000000",	-- 1685: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1686: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1687: 	jr	%ra
	-- o_param_r2.2658:
"00111000001000010000000000001001",	-- 1688: 	lw	%r1, [%r1 + 9]
"11001100000000100000000000000001",	-- 1689: 	lli	%r2, 1
"10000100001000100000100000000000",	-- 1690: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1691: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1692: 	jr	%ra
	-- o_param_r3.2660:
"00111000001000010000000000001001",	-- 1693: 	lw	%r1, [%r1 + 9]
"11001100000000100000000000000010",	-- 1694: 	lli	%r2, 2
"10000100001000100000100000000000",	-- 1695: 	add	%r1, %r1, %r2
"10010000001000000000000000000000",	-- 1696: 	lf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1697: 	jr	%ra
	-- o_param_ctbl.2662:
"00111000001000010000000000001010",	-- 1698: 	lw	%r1, [%r1 + 10]
"01001111111000000000000000000000",	-- 1699: 	jr	%ra
	-- p_rgb.2664:
"00111000001000010000000000000000",	-- 1700: 	lw	%r1, [%r1 + 0]
"01001111111000000000000000000000",	-- 1701: 	jr	%ra
	-- p_intersection_points.2666:
"00111000001000010000000000000001",	-- 1702: 	lw	%r1, [%r1 + 1]
"01001111111000000000000000000000",	-- 1703: 	jr	%ra
	-- p_surface_ids.2668:
"00111000001000010000000000000010",	-- 1704: 	lw	%r1, [%r1 + 2]
"01001111111000000000000000000000",	-- 1705: 	jr	%ra
	-- p_calc_diffuse.2670:
"00111000001000010000000000000011",	-- 1706: 	lw	%r1, [%r1 + 3]
"01001111111000000000000000000000",	-- 1707: 	jr	%ra
	-- p_energy.2672:
"00111000001000010000000000000100",	-- 1708: 	lw	%r1, [%r1 + 4]
"01001111111000000000000000000000",	-- 1709: 	jr	%ra
	-- p_received_ray_20percent.2674:
"00111000001000010000000000000101",	-- 1710: 	lw	%r1, [%r1 + 5]
"01001111111000000000000000000000",	-- 1711: 	jr	%ra
	-- p_group_id.2676:
"00111000001000010000000000000110",	-- 1712: 	lw	%r1, [%r1 + 6]
"11001100000000100000000000000000",	-- 1713: 	lli	%r2, 0
"10000100001000100000100000000000",	-- 1714: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 1715: 	lw	%r1, [%r1 + 0]
"01001111111000000000000000000000",	-- 1716: 	jr	%ra
	-- p_set_group_id.2678:
"00111000001000010000000000000110",	-- 1717: 	lw	%r1, [%r1 + 6]
"11001100000000110000000000000000",	-- 1718: 	lli	%r3, 0
"10000100001000110000100000000000",	-- 1719: 	add	%r1, %r1, %r3
"00111100010000010000000000000000",	-- 1720: 	sw	%r2, [%r1 + 0]
"01001111111000000000000000000000",	-- 1721: 	jr	%ra
	-- p_nvectors.2681:
"00111000001000010000000000000111",	-- 1722: 	lw	%r1, [%r1 + 7]
"01001111111000000000000000000000",	-- 1723: 	jr	%ra
	-- d_vec.2683:
"00111000001000010000000000000000",	-- 1724: 	lw	%r1, [%r1 + 0]
"01001111111000000000000000000000",	-- 1725: 	jr	%ra
	-- d_const.2685:
"00111000001000010000000000000001",	-- 1726: 	lw	%r1, [%r1 + 1]
"01001111111000000000000000000000",	-- 1727: 	jr	%ra
	-- r_surface_id.2687:
"00111000001000010000000000000000",	-- 1728: 	lw	%r1, [%r1 + 0]
"01001111111000000000000000000000",	-- 1729: 	jr	%ra
	-- r_dvec.2689:
"00111000001000010000000000000001",	-- 1730: 	lw	%r1, [%r1 + 1]
"01001111111000000000000000000000",	-- 1731: 	jr	%ra
	-- r_bright.2691:
"10010000001000000000000000000010",	-- 1732: 	lf	%f0, [%r1 + 2]
"01001111111000000000000000000000",	-- 1733: 	jr	%ra
	-- rad.2693:
"00010100000000011111100110011000",	-- 1734: 	llif	%f1, 0.017453
"00010000000000010011110010001110",	-- 1735: 	lhif	%f1, 0.017453
"11101000000000010000000000000000",	-- 1736: 	mulf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 1737: 	jr	%ra
	-- read_screen_settings.2695:
"00111011011000010000000000000101",	-- 1738: 	lw	%r1, [%r27 + 5]
"00111011011000100000000000000100",	-- 1739: 	lw	%r2, [%r27 + 4]
"00111011011000110000000000000011",	-- 1740: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 1741: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 1742: 	lw	%r5, [%r27 + 1]
"11001100000001100000000000000000",	-- 1743: 	lli	%r6, 0
"00111100001111100000000000000000",	-- 1744: 	sw	%r1, [%sp + 0]
"00111100011111100000000000000001",	-- 1745: 	sw	%r3, [%sp + 1]
"00111100100111100000000000000010",	-- 1746: 	sw	%r4, [%sp + 2]
"00111100010111100000000000000011",	-- 1747: 	sw	%r2, [%sp + 3]
"00111100110111100000000000000100",	-- 1748: 	sw	%r6, [%sp + 4]
"00111100101111100000000000000101",	-- 1749: 	sw	%r5, [%sp + 5]
"00111111111111100000000000000110",	-- 1750: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 1751: 	addi	%sp, %sp, 7
"01011000000000000010101001000001",	-- 1752: 	jal	yj_read_float
"10101011110111100000000000000111",	-- 1753: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 1754: 	lw	%ra, [%sp + 6]
"00111011110000010000000000000100",	-- 1755: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000101",	-- 1756: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 1757: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1758: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 1759: 	lli	%r1, 1
"00111100001111100000000000000110",	-- 1760: 	sw	%r1, [%sp + 6]
"00111111111111100000000000000111",	-- 1761: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 1762: 	addi	%sp, %sp, 8
"01011000000000000010101001000001",	-- 1763: 	jal	yj_read_float
"10101011110111100000000000001000",	-- 1764: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 1765: 	lw	%ra, [%sp + 7]
"00111011110000010000000000000110",	-- 1766: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000101",	-- 1767: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 1768: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1769: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 1770: 	lli	%r1, 2
"00111100001111100000000000000111",	-- 1771: 	sw	%r1, [%sp + 7]
"00111111111111100000000000001000",	-- 1772: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 1773: 	addi	%sp, %sp, 9
"01011000000000000010101001000001",	-- 1774: 	jal	yj_read_float
"10101011110111100000000000001001",	-- 1775: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 1776: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000111",	-- 1777: 	lw	%r1, [%sp + 7]
"00111011110000100000000000000101",	-- 1778: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 1779: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1780: 	sf	%f0, [%r1 + 0]
"00111111111111100000000000001000",	-- 1781: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 1782: 	addi	%sp, %sp, 9
"01011000000000000010101001000001",	-- 1783: 	jal	yj_read_float
"10101011110111100000000000001001",	-- 1784: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 1785: 	lw	%ra, [%sp + 8]
"00111111111111100000000000001000",	-- 1786: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 1787: 	addi	%sp, %sp, 9
"01011000000000000000011011000110",	-- 1788: 	jal	rad.2693
"10101011110111100000000000001001",	-- 1789: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 1790: 	lw	%ra, [%sp + 8]
"10110000000111100000000000001000",	-- 1791: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 1792: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 1793: 	addi	%sp, %sp, 10
"01011000000000000000010010011000",	-- 1794: 	jal	cos.2518
"10101011110111100000000000001010",	-- 1795: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 1796: 	lw	%ra, [%sp + 9]
"10010011110000010000000000001000",	-- 1797: 	lf	%f1, [%sp + 8]
"10110000000111100000000000001001",	-- 1798: 	sf	%f0, [%sp + 9]
"00001100001000000000000000000000",	-- 1799: 	movf	%f0, %f1
"00111111111111100000000000001010",	-- 1800: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 1801: 	addi	%sp, %sp, 11
"01011000000000000000010001011001",	-- 1802: 	jal	sin.2516
"10101011110111100000000000001011",	-- 1803: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 1804: 	lw	%ra, [%sp + 10]
"10110000000111100000000000001010",	-- 1805: 	sf	%f0, [%sp + 10]
"00111111111111100000000000001011",	-- 1806: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 1807: 	addi	%sp, %sp, 12
"01011000000000000010101001000001",	-- 1808: 	jal	yj_read_float
"10101011110111100000000000001100",	-- 1809: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 1810: 	lw	%ra, [%sp + 11]
"00111111111111100000000000001011",	-- 1811: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 1812: 	addi	%sp, %sp, 12
"01011000000000000000011011000110",	-- 1813: 	jal	rad.2693
"10101011110111100000000000001100",	-- 1814: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 1815: 	lw	%ra, [%sp + 11]
"10110000000111100000000000001011",	-- 1816: 	sf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 1817: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 1818: 	addi	%sp, %sp, 13
"01011000000000000000010010011000",	-- 1819: 	jal	cos.2518
"10101011110111100000000000001101",	-- 1820: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 1821: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001011",	-- 1822: 	lf	%f1, [%sp + 11]
"10110000000111100000000000001100",	-- 1823: 	sf	%f0, [%sp + 12]
"00001100001000000000000000000000",	-- 1824: 	movf	%f0, %f1
"00111111111111100000000000001101",	-- 1825: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 1826: 	addi	%sp, %sp, 14
"01011000000000000000010001011001",	-- 1827: 	jal	sin.2516
"10101011110111100000000000001110",	-- 1828: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 1829: 	lw	%ra, [%sp + 13]
"11001100000000010000000000000000",	-- 1830: 	lli	%r1, 0
"10010011110000010000000000001001",	-- 1831: 	lf	%f1, [%sp + 9]
"11101000001000000001000000000000",	-- 1832: 	mulf	%f2, %f1, %f0
"00010100000000110000000000000000",	-- 1833: 	llif	%f3, 200.000000
"00010000000000110100001101001000",	-- 1834: 	lhif	%f3, 200.000000
"11101000010000110001000000000000",	-- 1835: 	mulf	%f2, %f2, %f3
"00111011110000100000000000000011",	-- 1836: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 1837: 	add	%r1, %r2, %r1
"10110000010000010000000000000000",	-- 1838: 	sf	%f2, [%r1 + 0]
"11001100000000010000000000000001",	-- 1839: 	lli	%r1, 1
"00010100000000100000000000000000",	-- 1840: 	llif	%f2, -200.000000
"00010000000000101100001101001000",	-- 1841: 	lhif	%f2, -200.000000
"10010011110000110000000000001010",	-- 1842: 	lf	%f3, [%sp + 10]
"11101000011000100001000000000000",	-- 1843: 	mulf	%f2, %f3, %f2
"10000100010000010000100000000000",	-- 1844: 	add	%r1, %r2, %r1
"10110000010000010000000000000000",	-- 1845: 	sf	%f2, [%r1 + 0]
"11001100000000010000000000000010",	-- 1846: 	lli	%r1, 2
"10010011110000100000000000001100",	-- 1847: 	lf	%f2, [%sp + 12]
"11101000001000100010000000000000",	-- 1848: 	mulf	%f4, %f1, %f2
"00010100000001010000000000000000",	-- 1849: 	llif	%f5, 200.000000
"00010000000001010100001101001000",	-- 1850: 	lhif	%f5, 200.000000
"11101000100001010010000000000000",	-- 1851: 	mulf	%f4, %f4, %f5
"10000100010000010000100000000000",	-- 1852: 	add	%r1, %r2, %r1
"10110000100000010000000000000000",	-- 1853: 	sf	%f4, [%r1 + 0]
"11001100000000010000000000000000",	-- 1854: 	lli	%r1, 0
"00111011110000110000000000000010",	-- 1855: 	lw	%r3, [%sp + 2]
"10000100011000010000100000000000",	-- 1856: 	add	%r1, %r3, %r1
"10110000010000010000000000000000",	-- 1857: 	sf	%f2, [%r1 + 0]
"11001100000000010000000000000001",	-- 1858: 	lli	%r1, 1
"00010100000001000000000000000000",	-- 1859: 	llif	%f4, 0.000000
"00010000000001000000000000000000",	-- 1860: 	lhif	%f4, 0.000000
"10000100011000010000100000000000",	-- 1861: 	add	%r1, %r3, %r1
"10110000100000010000000000000000",	-- 1862: 	sf	%f4, [%r1 + 0]
"11001100000000010000000000000010",	-- 1863: 	lli	%r1, 2
"10110000000111100000000000001101",	-- 1864: 	sf	%f0, [%sp + 13]
"00111100001111100000000000001110",	-- 1865: 	sw	%r1, [%sp + 14]
"00111111111111100000000000001111",	-- 1866: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 1867: 	addi	%sp, %sp, 16
"01011000000000000010101001010001",	-- 1868: 	jal	yj_fneg
"10101011110111100000000000010000",	-- 1869: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 1870: 	lw	%ra, [%sp + 15]
"00111011110000010000000000001110",	-- 1871: 	lw	%r1, [%sp + 14]
"00111011110000100000000000000010",	-- 1872: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 1873: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1874: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 1875: 	lli	%r1, 0
"10010011110000000000000000001010",	-- 1876: 	lf	%f0, [%sp + 10]
"00111100001111100000000000001111",	-- 1877: 	sw	%r1, [%sp + 15]
"00111111111111100000000000010000",	-- 1878: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 1879: 	addi	%sp, %sp, 17
"01011000000000000010101001010001",	-- 1880: 	jal	yj_fneg
"10101011110111100000000000010001",	-- 1881: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 1882: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001101",	-- 1883: 	lf	%f1, [%sp + 13]
"11101000000000010000000000000000",	-- 1884: 	mulf	%f0, %f0, %f1
"00111011110000010000000000001111",	-- 1885: 	lw	%r1, [%sp + 15]
"00111011110000100000000000000001",	-- 1886: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 1887: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1888: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 1889: 	lli	%r1, 1
"10010011110000000000000000001001",	-- 1890: 	lf	%f0, [%sp + 9]
"00111100001111100000000000010000",	-- 1891: 	sw	%r1, [%sp + 16]
"00111111111111100000000000010001",	-- 1892: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 1893: 	addi	%sp, %sp, 18
"01011000000000000010101001010001",	-- 1894: 	jal	yj_fneg
"10101011110111100000000000010010",	-- 1895: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 1896: 	lw	%ra, [%sp + 17]
"00111011110000010000000000010000",	-- 1897: 	lw	%r1, [%sp + 16]
"00111011110000100000000000000001",	-- 1898: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 1899: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1900: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 1901: 	lli	%r1, 2
"10010011110000000000000000001010",	-- 1902: 	lf	%f0, [%sp + 10]
"00111100001111100000000000010001",	-- 1903: 	sw	%r1, [%sp + 17]
"00111111111111100000000000010010",	-- 1904: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 1905: 	addi	%sp, %sp, 19
"01011000000000000010101001010001",	-- 1906: 	jal	yj_fneg
"10101011110111100000000000010011",	-- 1907: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 1908: 	lw	%ra, [%sp + 18]
"10010011110000010000000000001100",	-- 1909: 	lf	%f1, [%sp + 12]
"11101000000000010000000000000000",	-- 1910: 	mulf	%f0, %f0, %f1
"00111011110000010000000000010001",	-- 1911: 	lw	%r1, [%sp + 17]
"00111011110000100000000000000001",	-- 1912: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 1913: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1914: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 1915: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 1916: 	lli	%r2, 0
"00111011110000110000000000000101",	-- 1917: 	lw	%r3, [%sp + 5]
"10000100011000100001000000000000",	-- 1918: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 1919: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000000",	-- 1920: 	lli	%r2, 0
"00111011110001000000000000000011",	-- 1921: 	lw	%r4, [%sp + 3]
"10000100100000100001000000000000",	-- 1922: 	add	%r2, %r4, %r2
"10010000010000010000000000000000",	-- 1923: 	lf	%f1, [%r2 + 0]
"11100100000000010000000000000000",	-- 1924: 	subf	%f0, %f0, %f1
"00111011110000100000000000000000",	-- 1925: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 1926: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1927: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 1928: 	lli	%r1, 1
"11001100000001010000000000000001",	-- 1929: 	lli	%r5, 1
"10000100011001010010100000000000",	-- 1930: 	add	%r5, %r3, %r5
"10010000101000000000000000000000",	-- 1931: 	lf	%f0, [%r5 + 0]
"11001100000001010000000000000001",	-- 1932: 	lli	%r5, 1
"10000100100001010010100000000000",	-- 1933: 	add	%r5, %r4, %r5
"10010000101000010000000000000000",	-- 1934: 	lf	%f1, [%r5 + 0]
"11100100000000010000000000000000",	-- 1935: 	subf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 1936: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1937: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 1938: 	lli	%r1, 2
"11001100000001010000000000000010",	-- 1939: 	lli	%r5, 2
"10000100011001010001100000000000",	-- 1940: 	add	%r3, %r3, %r5
"10010000011000000000000000000000",	-- 1941: 	lf	%f0, [%r3 + 0]
"11001100000000110000000000000010",	-- 1942: 	lli	%r3, 2
"10000100100000110001100000000000",	-- 1943: 	add	%r3, %r4, %r3
"10010000011000010000000000000000",	-- 1944: 	lf	%f1, [%r3 + 0]
"11100100000000010000000000000000",	-- 1945: 	subf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 1946: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1947: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 1948: 	jr	%ra
	-- read_light.2697:
"00111011011000010000000000000010",	-- 1949: 	lw	%r1, [%r27 + 2]
"00111011011000100000000000000001",	-- 1950: 	lw	%r2, [%r27 + 1]
"00111100010111100000000000000000",	-- 1951: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 1952: 	sw	%r1, [%sp + 1]
"00111111111111100000000000000010",	-- 1953: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1954: 	addi	%sp, %sp, 3
"01011000000000000010101000110100",	-- 1955: 	jal	yj_read_int
"10101011110111100000000000000011",	-- 1956: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1957: 	lw	%ra, [%sp + 2]
"00111111111111100000000000000010",	-- 1958: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1959: 	addi	%sp, %sp, 3
"01011000000000000010101001000001",	-- 1960: 	jal	yj_read_float
"10101011110111100000000000000011",	-- 1961: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1962: 	lw	%ra, [%sp + 2]
"00111111111111100000000000000010",	-- 1963: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 1964: 	addi	%sp, %sp, 3
"01011000000000000000011011000110",	-- 1965: 	jal	rad.2693
"10101011110111100000000000000011",	-- 1966: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 1967: 	lw	%ra, [%sp + 2]
"10110000000111100000000000000010",	-- 1968: 	sf	%f0, [%sp + 2]
"00111111111111100000000000000011",	-- 1969: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 1970: 	addi	%sp, %sp, 4
"01011000000000000000010001011001",	-- 1971: 	jal	sin.2516
"10101011110111100000000000000100",	-- 1972: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 1973: 	lw	%ra, [%sp + 3]
"11001100000000010000000000000001",	-- 1974: 	lli	%r1, 1
"00111100001111100000000000000011",	-- 1975: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 1976: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 1977: 	addi	%sp, %sp, 5
"01011000000000000010101001010001",	-- 1978: 	jal	yj_fneg
"10101011110111100000000000000101",	-- 1979: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 1980: 	lw	%ra, [%sp + 4]
"00111011110000010000000000000011",	-- 1981: 	lw	%r1, [%sp + 3]
"00111011110000100000000000000001",	-- 1982: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 1983: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 1984: 	sf	%f0, [%r1 + 0]
"00111111111111100000000000000100",	-- 1985: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 1986: 	addi	%sp, %sp, 5
"01011000000000000010101001000001",	-- 1987: 	jal	yj_read_float
"10101011110111100000000000000101",	-- 1988: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 1989: 	lw	%ra, [%sp + 4]
"00111111111111100000000000000100",	-- 1990: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 1991: 	addi	%sp, %sp, 5
"01011000000000000000011011000110",	-- 1992: 	jal	rad.2693
"10101011110111100000000000000101",	-- 1993: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 1994: 	lw	%ra, [%sp + 4]
"10010011110000010000000000000010",	-- 1995: 	lf	%f1, [%sp + 2]
"10110000000111100000000000000100",	-- 1996: 	sf	%f0, [%sp + 4]
"00001100001000000000000000000000",	-- 1997: 	movf	%f0, %f1
"00111111111111100000000000000101",	-- 1998: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 1999: 	addi	%sp, %sp, 6
"01011000000000000000010010011000",	-- 2000: 	jal	cos.2518
"10101011110111100000000000000110",	-- 2001: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 2002: 	lw	%ra, [%sp + 5]
"10010011110000010000000000000100",	-- 2003: 	lf	%f1, [%sp + 4]
"10110000000111100000000000000101",	-- 2004: 	sf	%f0, [%sp + 5]
"00001100001000000000000000000000",	-- 2005: 	movf	%f0, %f1
"00111111111111100000000000000110",	-- 2006: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 2007: 	addi	%sp, %sp, 7
"01011000000000000000010001011001",	-- 2008: 	jal	sin.2516
"10101011110111100000000000000111",	-- 2009: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 2010: 	lw	%ra, [%sp + 6]
"11001100000000010000000000000000",	-- 2011: 	lli	%r1, 0
"10010011110000010000000000000101",	-- 2012: 	lf	%f1, [%sp + 5]
"11101000001000000000000000000000",	-- 2013: 	mulf	%f0, %f1, %f0
"00111011110000100000000000000001",	-- 2014: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2015: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2016: 	sf	%f0, [%r1 + 0]
"10010011110000000000000000000100",	-- 2017: 	lf	%f0, [%sp + 4]
"00111111111111100000000000000110",	-- 2018: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 2019: 	addi	%sp, %sp, 7
"01011000000000000000010010011000",	-- 2020: 	jal	cos.2518
"10101011110111100000000000000111",	-- 2021: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 2022: 	lw	%ra, [%sp + 6]
"11001100000000010000000000000010",	-- 2023: 	lli	%r1, 2
"10010011110000010000000000000101",	-- 2024: 	lf	%f1, [%sp + 5]
"11101000001000000000000000000000",	-- 2025: 	mulf	%f0, %f1, %f0
"00111011110000100000000000000001",	-- 2026: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2027: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2028: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 2029: 	lli	%r1, 0
"00111100001111100000000000000110",	-- 2030: 	sw	%r1, [%sp + 6]
"00111111111111100000000000000111",	-- 2031: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 2032: 	addi	%sp, %sp, 8
"01011000000000000010101001000001",	-- 2033: 	jal	yj_read_float
"10101011110111100000000000001000",	-- 2034: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 2035: 	lw	%ra, [%sp + 7]
"00111011110000010000000000000110",	-- 2036: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000000",	-- 2037: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 2038: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2039: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 2040: 	jr	%ra
	-- rotate_quadratic_matrix.2699:
"11001100000000110000000000000000",	-- 2041: 	lli	%r3, 0
"10000100010000110001100000000000",	-- 2042: 	add	%r3, %r2, %r3
"10010000011000000000000000000000",	-- 2043: 	lf	%f0, [%r3 + 0]
"00111100001111100000000000000000",	-- 2044: 	sw	%r1, [%sp + 0]
"00111100010111100000000000000001",	-- 2045: 	sw	%r2, [%sp + 1]
"00111111111111100000000000000010",	-- 2046: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 2047: 	addi	%sp, %sp, 3
"01011000000000000000010010011000",	-- 2048: 	jal	cos.2518
"10101011110111100000000000000011",	-- 2049: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 2050: 	lw	%ra, [%sp + 2]
"11001100000000010000000000000000",	-- 2051: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 2052: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2053: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 2054: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000010",	-- 2055: 	sf	%f0, [%sp + 2]
"00001100001000000000000000000000",	-- 2056: 	movf	%f0, %f1
"00111111111111100000000000000011",	-- 2057: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 2058: 	addi	%sp, %sp, 4
"01011000000000000000010001011001",	-- 2059: 	jal	sin.2516
"10101011110111100000000000000100",	-- 2060: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 2061: 	lw	%ra, [%sp + 3]
"11001100000000010000000000000001",	-- 2062: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 2063: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2064: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 2065: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000011",	-- 2066: 	sf	%f0, [%sp + 3]
"00001100001000000000000000000000",	-- 2067: 	movf	%f0, %f1
"00111111111111100000000000000100",	-- 2068: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 2069: 	addi	%sp, %sp, 5
"01011000000000000000010010011000",	-- 2070: 	jal	cos.2518
"10101011110111100000000000000101",	-- 2071: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 2072: 	lw	%ra, [%sp + 4]
"11001100000000010000000000000001",	-- 2073: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 2074: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2075: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 2076: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000100",	-- 2077: 	sf	%f0, [%sp + 4]
"00001100001000000000000000000000",	-- 2078: 	movf	%f0, %f1
"00111111111111100000000000000101",	-- 2079: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 2080: 	addi	%sp, %sp, 6
"01011000000000000000010001011001",	-- 2081: 	jal	sin.2516
"10101011110111100000000000000110",	-- 2082: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 2083: 	lw	%ra, [%sp + 5]
"11001100000000010000000000000010",	-- 2084: 	lli	%r1, 2
"00111011110000100000000000000001",	-- 2085: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2086: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 2087: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000101",	-- 2088: 	sf	%f0, [%sp + 5]
"00001100001000000000000000000000",	-- 2089: 	movf	%f0, %f1
"00111111111111100000000000000110",	-- 2090: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 2091: 	addi	%sp, %sp, 7
"01011000000000000000010010011000",	-- 2092: 	jal	cos.2518
"10101011110111100000000000000111",	-- 2093: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 2094: 	lw	%ra, [%sp + 6]
"11001100000000010000000000000010",	-- 2095: 	lli	%r1, 2
"00111011110000100000000000000001",	-- 2096: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2097: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 2098: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000110",	-- 2099: 	sf	%f0, [%sp + 6]
"00001100001000000000000000000000",	-- 2100: 	movf	%f0, %f1
"00111111111111100000000000000111",	-- 2101: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 2102: 	addi	%sp, %sp, 8
"01011000000000000000010001011001",	-- 2103: 	jal	sin.2516
"10101011110111100000000000001000",	-- 2104: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 2105: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000110",	-- 2106: 	lf	%f1, [%sp + 6]
"10010011110000100000000000000100",	-- 2107: 	lf	%f2, [%sp + 4]
"11101000010000010001100000000000",	-- 2108: 	mulf	%f3, %f2, %f1
"10010011110001000000000000000101",	-- 2109: 	lf	%f4, [%sp + 5]
"10010011110001010000000000000011",	-- 2110: 	lf	%f5, [%sp + 3]
"11101000101001000011000000000000",	-- 2111: 	mulf	%f6, %f5, %f4
"11101000110000010011000000000000",	-- 2112: 	mulf	%f6, %f6, %f1
"10010011110001110000000000000010",	-- 2113: 	lf	%f7, [%sp + 2]
"11101000111000000100000000000000",	-- 2114: 	mulf	%f8, %f7, %f0
"11100100110010000011000000000000",	-- 2115: 	subf	%f6, %f6, %f8
"11101000111001000100000000000000",	-- 2116: 	mulf	%f8, %f7, %f4
"11101001000000010100000000000000",	-- 2117: 	mulf	%f8, %f8, %f1
"11101000101000000100100000000000",	-- 2118: 	mulf	%f9, %f5, %f0
"11100001000010010100000000000000",	-- 2119: 	addf	%f8, %f8, %f9
"11101000010000000100100000000000",	-- 2120: 	mulf	%f9, %f2, %f0
"11101000101001000101000000000000",	-- 2121: 	mulf	%f10, %f5, %f4
"11101001010000000101000000000000",	-- 2122: 	mulf	%f10, %f10, %f0
"11101000111000010101100000000000",	-- 2123: 	mulf	%f11, %f7, %f1
"11100001010010110101000000000000",	-- 2124: 	addf	%f10, %f10, %f11
"11101000111001000101100000000000",	-- 2125: 	mulf	%f11, %f7, %f4
"11101001011000000000000000000000",	-- 2126: 	mulf	%f0, %f11, %f0
"11101000101000010000100000000000",	-- 2127: 	mulf	%f1, %f5, %f1
"11100100000000010000000000000000",	-- 2128: 	subf	%f0, %f0, %f1
"10110000000111100000000000000111",	-- 2129: 	sf	%f0, [%sp + 7]
"10110001000111100000000000001000",	-- 2130: 	sf	%f8, [%sp + 8]
"10110001010111100000000000001001",	-- 2131: 	sf	%f10, [%sp + 9]
"10110000110111100000000000001010",	-- 2132: 	sf	%f6, [%sp + 10]
"10110001001111100000000000001011",	-- 2133: 	sf	%f9, [%sp + 11]
"10110000011111100000000000001100",	-- 2134: 	sf	%f3, [%sp + 12]
"00001100100000000000000000000000",	-- 2135: 	movf	%f0, %f4
"00111111111111100000000000001101",	-- 2136: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 2137: 	addi	%sp, %sp, 14
"01011000000000000010101001010001",	-- 2138: 	jal	yj_fneg
"10101011110111100000000000001110",	-- 2139: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 2140: 	lw	%ra, [%sp + 13]
"10010011110000010000000000000100",	-- 2141: 	lf	%f1, [%sp + 4]
"10010011110000100000000000000011",	-- 2142: 	lf	%f2, [%sp + 3]
"11101000010000010001000000000000",	-- 2143: 	mulf	%f2, %f2, %f1
"10010011110000110000000000000010",	-- 2144: 	lf	%f3, [%sp + 2]
"11101000011000010000100000000000",	-- 2145: 	mulf	%f1, %f3, %f1
"11001100000000010000000000000000",	-- 2146: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 2147: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 2148: 	add	%r1, %r2, %r1
"10010000001000110000000000000000",	-- 2149: 	lf	%f3, [%r1 + 0]
"11001100000000010000000000000001",	-- 2150: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 2151: 	add	%r1, %r2, %r1
"10010000001001000000000000000000",	-- 2152: 	lf	%f4, [%r1 + 0]
"11001100000000010000000000000010",	-- 2153: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 2154: 	add	%r1, %r2, %r1
"10010000001001010000000000000000",	-- 2155: 	lf	%f5, [%r1 + 0]
"11001100000000010000000000000000",	-- 2156: 	lli	%r1, 0
"10010011110001100000000000001100",	-- 2157: 	lf	%f6, [%sp + 12]
"10110000001111100000000000001101",	-- 2158: 	sf	%f1, [%sp + 13]
"10110000010111100000000000001110",	-- 2159: 	sf	%f2, [%sp + 14]
"00111100001111100000000000001111",	-- 2160: 	sw	%r1, [%sp + 15]
"10110000101111100000000000010000",	-- 2161: 	sf	%f5, [%sp + 16]
"10110000000111100000000000010001",	-- 2162: 	sf	%f0, [%sp + 17]
"10110000100111100000000000010010",	-- 2163: 	sf	%f4, [%sp + 18]
"10110000011111100000000000010011",	-- 2164: 	sf	%f3, [%sp + 19]
"00001100110000000000000000000000",	-- 2165: 	movf	%f0, %f6
"00111111111111100000000000010100",	-- 2166: 	sw	%ra, [%sp + 20]
"10100111110111100000000000010101",	-- 2167: 	addi	%sp, %sp, 21
"01011000000000000000010011110001",	-- 2168: 	jal	fsqr.2530
"10101011110111100000000000010101",	-- 2169: 	subi	%sp, %sp, 21
"00111011110111110000000000010100",	-- 2170: 	lw	%ra, [%sp + 20]
"10010011110000010000000000010011",	-- 2171: 	lf	%f1, [%sp + 19]
"11101000001000000000000000000000",	-- 2172: 	mulf	%f0, %f1, %f0
"10010011110000100000000000001011",	-- 2173: 	lf	%f2, [%sp + 11]
"10110000000111100000000000010100",	-- 2174: 	sf	%f0, [%sp + 20]
"00001100010000000000000000000000",	-- 2175: 	movf	%f0, %f2
"00111111111111100000000000010101",	-- 2176: 	sw	%ra, [%sp + 21]
"10100111110111100000000000010110",	-- 2177: 	addi	%sp, %sp, 22
"01011000000000000000010011110001",	-- 2178: 	jal	fsqr.2530
"10101011110111100000000000010110",	-- 2179: 	subi	%sp, %sp, 22
"00111011110111110000000000010101",	-- 2180: 	lw	%ra, [%sp + 21]
"10010011110000010000000000010010",	-- 2181: 	lf	%f1, [%sp + 18]
"11101000001000000000000000000000",	-- 2182: 	mulf	%f0, %f1, %f0
"10010011110000100000000000010100",	-- 2183: 	lf	%f2, [%sp + 20]
"11100000010000000000000000000000",	-- 2184: 	addf	%f0, %f2, %f0
"10010011110000100000000000010001",	-- 2185: 	lf	%f2, [%sp + 17]
"10110000000111100000000000010101",	-- 2186: 	sf	%f0, [%sp + 21]
"00001100010000000000000000000000",	-- 2187: 	movf	%f0, %f2
"00111111111111100000000000010110",	-- 2188: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 2189: 	addi	%sp, %sp, 23
"01011000000000000000010011110001",	-- 2190: 	jal	fsqr.2530
"10101011110111100000000000010111",	-- 2191: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 2192: 	lw	%ra, [%sp + 22]
"10010011110000010000000000010000",	-- 2193: 	lf	%f1, [%sp + 16]
"11101000001000000000000000000000",	-- 2194: 	mulf	%f0, %f1, %f0
"10010011110000100000000000010101",	-- 2195: 	lf	%f2, [%sp + 21]
"11100000010000000000000000000000",	-- 2196: 	addf	%f0, %f2, %f0
"00111011110000010000000000001111",	-- 2197: 	lw	%r1, [%sp + 15]
"00111011110000100000000000000000",	-- 2198: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 2199: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2200: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2201: 	lli	%r1, 1
"10010011110000000000000000001010",	-- 2202: 	lf	%f0, [%sp + 10]
"00111100001111100000000000010110",	-- 2203: 	sw	%r1, [%sp + 22]
"00111111111111100000000000010111",	-- 2204: 	sw	%ra, [%sp + 23]
"10100111110111100000000000011000",	-- 2205: 	addi	%sp, %sp, 24
"01011000000000000000010011110001",	-- 2206: 	jal	fsqr.2530
"10101011110111100000000000011000",	-- 2207: 	subi	%sp, %sp, 24
"00111011110111110000000000010111",	-- 2208: 	lw	%ra, [%sp + 23]
"10010011110000010000000000010011",	-- 2209: 	lf	%f1, [%sp + 19]
"11101000001000000000000000000000",	-- 2210: 	mulf	%f0, %f1, %f0
"10010011110000100000000000001001",	-- 2211: 	lf	%f2, [%sp + 9]
"10110000000111100000000000010111",	-- 2212: 	sf	%f0, [%sp + 23]
"00001100010000000000000000000000",	-- 2213: 	movf	%f0, %f2
"00111111111111100000000000011000",	-- 2214: 	sw	%ra, [%sp + 24]
"10100111110111100000000000011001",	-- 2215: 	addi	%sp, %sp, 25
"01011000000000000000010011110001",	-- 2216: 	jal	fsqr.2530
"10101011110111100000000000011001",	-- 2217: 	subi	%sp, %sp, 25
"00111011110111110000000000011000",	-- 2218: 	lw	%ra, [%sp + 24]
"10010011110000010000000000010010",	-- 2219: 	lf	%f1, [%sp + 18]
"11101000001000000000000000000000",	-- 2220: 	mulf	%f0, %f1, %f0
"10010011110000100000000000010111",	-- 2221: 	lf	%f2, [%sp + 23]
"11100000010000000000000000000000",	-- 2222: 	addf	%f0, %f2, %f0
"10010011110000100000000000001110",	-- 2223: 	lf	%f2, [%sp + 14]
"10110000000111100000000000011000",	-- 2224: 	sf	%f0, [%sp + 24]
"00001100010000000000000000000000",	-- 2225: 	movf	%f0, %f2
"00111111111111100000000000011001",	-- 2226: 	sw	%ra, [%sp + 25]
"10100111110111100000000000011010",	-- 2227: 	addi	%sp, %sp, 26
"01011000000000000000010011110001",	-- 2228: 	jal	fsqr.2530
"10101011110111100000000000011010",	-- 2229: 	subi	%sp, %sp, 26
"00111011110111110000000000011001",	-- 2230: 	lw	%ra, [%sp + 25]
"10010011110000010000000000010000",	-- 2231: 	lf	%f1, [%sp + 16]
"11101000001000000000000000000000",	-- 2232: 	mulf	%f0, %f1, %f0
"10010011110000100000000000011000",	-- 2233: 	lf	%f2, [%sp + 24]
"11100000010000000000000000000000",	-- 2234: 	addf	%f0, %f2, %f0
"00111011110000010000000000010110",	-- 2235: 	lw	%r1, [%sp + 22]
"00111011110000100000000000000000",	-- 2236: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 2237: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2238: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2239: 	lli	%r1, 2
"10010011110000000000000000001000",	-- 2240: 	lf	%f0, [%sp + 8]
"00111100001111100000000000011001",	-- 2241: 	sw	%r1, [%sp + 25]
"00111111111111100000000000011010",	-- 2242: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 2243: 	addi	%sp, %sp, 27
"01011000000000000000010011110001",	-- 2244: 	jal	fsqr.2530
"10101011110111100000000000011011",	-- 2245: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 2246: 	lw	%ra, [%sp + 26]
"10010011110000010000000000010011",	-- 2247: 	lf	%f1, [%sp + 19]
"11101000001000000000000000000000",	-- 2248: 	mulf	%f0, %f1, %f0
"10010011110000100000000000000111",	-- 2249: 	lf	%f2, [%sp + 7]
"10110000000111100000000000011010",	-- 2250: 	sf	%f0, [%sp + 26]
"00001100010000000000000000000000",	-- 2251: 	movf	%f0, %f2
"00111111111111100000000000011011",	-- 2252: 	sw	%ra, [%sp + 27]
"10100111110111100000000000011100",	-- 2253: 	addi	%sp, %sp, 28
"01011000000000000000010011110001",	-- 2254: 	jal	fsqr.2530
"10101011110111100000000000011100",	-- 2255: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 2256: 	lw	%ra, [%sp + 27]
"10010011110000010000000000010010",	-- 2257: 	lf	%f1, [%sp + 18]
"11101000001000000000000000000000",	-- 2258: 	mulf	%f0, %f1, %f0
"10010011110000100000000000011010",	-- 2259: 	lf	%f2, [%sp + 26]
"11100000010000000000000000000000",	-- 2260: 	addf	%f0, %f2, %f0
"10010011110000100000000000001101",	-- 2261: 	lf	%f2, [%sp + 13]
"10110000000111100000000000011011",	-- 2262: 	sf	%f0, [%sp + 27]
"00001100010000000000000000000000",	-- 2263: 	movf	%f0, %f2
"00111111111111100000000000011100",	-- 2264: 	sw	%ra, [%sp + 28]
"10100111110111100000000000011101",	-- 2265: 	addi	%sp, %sp, 29
"01011000000000000000010011110001",	-- 2266: 	jal	fsqr.2530
"10101011110111100000000000011101",	-- 2267: 	subi	%sp, %sp, 29
"00111011110111110000000000011100",	-- 2268: 	lw	%ra, [%sp + 28]
"10010011110000010000000000010000",	-- 2269: 	lf	%f1, [%sp + 16]
"11101000001000000000000000000000",	-- 2270: 	mulf	%f0, %f1, %f0
"10010011110000100000000000011011",	-- 2271: 	lf	%f2, [%sp + 27]
"11100000010000000000000000000000",	-- 2272: 	addf	%f0, %f2, %f0
"00111011110000010000000000011001",	-- 2273: 	lw	%r1, [%sp + 25]
"00111011110000100000000000000000",	-- 2274: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 2275: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2276: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 2277: 	lli	%r1, 0
"00010100000000000000000000000000",	-- 2278: 	llif	%f0, 2.000000
"00010000000000000100000000000000",	-- 2279: 	lhif	%f0, 2.000000
"10010011110000100000000000001010",	-- 2280: 	lf	%f2, [%sp + 10]
"10010011110000110000000000010011",	-- 2281: 	lf	%f3, [%sp + 19]
"11101000011000100010000000000000",	-- 2282: 	mulf	%f4, %f3, %f2
"10010011110001010000000000001000",	-- 2283: 	lf	%f5, [%sp + 8]
"11101000100001010010000000000000",	-- 2284: 	mulf	%f4, %f4, %f5
"10010011110001100000000000001001",	-- 2285: 	lf	%f6, [%sp + 9]
"10010011110001110000000000010010",	-- 2286: 	lf	%f7, [%sp + 18]
"11101000111001100100000000000000",	-- 2287: 	mulf	%f8, %f7, %f6
"10010011110010010000000000000111",	-- 2288: 	lf	%f9, [%sp + 7]
"11101001000010010100000000000000",	-- 2289: 	mulf	%f8, %f8, %f9
"11100000100010000010000000000000",	-- 2290: 	addf	%f4, %f4, %f8
"10010011110010000000000000001110",	-- 2291: 	lf	%f8, [%sp + 14]
"11101000001010000101000000000000",	-- 2292: 	mulf	%f10, %f1, %f8
"10010011110010110000000000001101",	-- 2293: 	lf	%f11, [%sp + 13]
"11101001010010110101000000000000",	-- 2294: 	mulf	%f10, %f10, %f11
"11100000100010100010000000000000",	-- 2295: 	addf	%f4, %f4, %f10
"11101000000001000000000000000000",	-- 2296: 	mulf	%f0, %f0, %f4
"00111011110000100000000000000001",	-- 2297: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2298: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2299: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2300: 	lli	%r1, 1
"00010100000000000000000000000000",	-- 2301: 	llif	%f0, 2.000000
"00010000000000000100000000000000",	-- 2302: 	lhif	%f0, 2.000000
"10010011110001000000000000001100",	-- 2303: 	lf	%f4, [%sp + 12]
"11101000011001000101000000000000",	-- 2304: 	mulf	%f10, %f3, %f4
"11101001010001010010100000000000",	-- 2305: 	mulf	%f5, %f10, %f5
"10010011110010100000000000001011",	-- 2306: 	lf	%f10, [%sp + 11]
"11101000111010100110000000000000",	-- 2307: 	mulf	%f12, %f7, %f10
"11101001100010010100100000000000",	-- 2308: 	mulf	%f9, %f12, %f9
"11100000101010010010100000000000",	-- 2309: 	addf	%f5, %f5, %f9
"10010011110010010000000000010001",	-- 2310: 	lf	%f9, [%sp + 17]
"11101000001010010110000000000000",	-- 2311: 	mulf	%f12, %f1, %f9
"11101001100010110101100000000000",	-- 2312: 	mulf	%f11, %f12, %f11
"11100000101010110010100000000000",	-- 2313: 	addf	%f5, %f5, %f11
"11101000000001010000000000000000",	-- 2314: 	mulf	%f0, %f0, %f5
"10000100010000010000100000000000",	-- 2315: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2316: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2317: 	lli	%r1, 2
"00010100000000000000000000000000",	-- 2318: 	llif	%f0, 2.000000
"00010000000000000100000000000000",	-- 2319: 	lhif	%f0, 2.000000
"11101000011001000001100000000000",	-- 2320: 	mulf	%f3, %f3, %f4
"11101000011000100001000000000000",	-- 2321: 	mulf	%f2, %f3, %f2
"11101000111010100001100000000000",	-- 2322: 	mulf	%f3, %f7, %f10
"11101000011001100001100000000000",	-- 2323: 	mulf	%f3, %f3, %f6
"11100000010000110001000000000000",	-- 2324: 	addf	%f2, %f2, %f3
"11101000001010010000100000000000",	-- 2325: 	mulf	%f1, %f1, %f9
"11101000001010000000100000000000",	-- 2326: 	mulf	%f1, %f1, %f8
"11100000010000010000100000000000",	-- 2327: 	addf	%f1, %f2, %f1
"11101000000000010000000000000000",	-- 2328: 	mulf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 2329: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2330: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 2331: 	jr	%ra
	-- read_nth_object.2702:
"00111011011000100000000000000001",	-- 2332: 	lw	%r2, [%r27 + 1]
"00111100001111100000000000000000",	-- 2333: 	sw	%r1, [%sp + 0]
"00111100010111100000000000000001",	-- 2334: 	sw	%r2, [%sp + 1]
"00111111111111100000000000000010",	-- 2335: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 2336: 	addi	%sp, %sp, 3
"01011000000000000010101000110100",	-- 2337: 	jal	yj_read_int
"10101011110111100000000000000011",	-- 2338: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 2339: 	lw	%ra, [%sp + 2]
"11001100000000101111111111111111",	-- 2340: 	lli	%r2, -1
"11001000000000101111111111111111",	-- 2341: 	lhi	%r2, -1
"00101000001000100000000000000011",	-- 2342: 	bneq	%r1, %r2, bneq_else.8961
"11001100000000010000000000000000",	-- 2343: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 2344: 	jr	%ra
	-- bneq_else.8961:
"00111100001111100000000000000010",	-- 2345: 	sw	%r1, [%sp + 2]
"00111111111111100000000000000011",	-- 2346: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 2347: 	addi	%sp, %sp, 4
"01011000000000000010101000110100",	-- 2348: 	jal	yj_read_int
"10101011110111100000000000000100",	-- 2349: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 2350: 	lw	%ra, [%sp + 3]
"00111100001111100000000000000011",	-- 2351: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 2352: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 2353: 	addi	%sp, %sp, 5
"01011000000000000010101000110100",	-- 2354: 	jal	yj_read_int
"10101011110111100000000000000101",	-- 2355: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 2356: 	lw	%ra, [%sp + 4]
"00111100001111100000000000000100",	-- 2357: 	sw	%r1, [%sp + 4]
"00111111111111100000000000000101",	-- 2358: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 2359: 	addi	%sp, %sp, 6
"01011000000000000010101000110100",	-- 2360: 	jal	yj_read_int
"10101011110111100000000000000110",	-- 2361: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 2362: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000011",	-- 2363: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 2364: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2365: 	lhif	%f0, 0.000000
"00111100001111100000000000000101",	-- 2366: 	sw	%r1, [%sp + 5]
"10000100000000100000100000000000",	-- 2367: 	add	%r1, %r0, %r2
"00111111111111100000000000000110",	-- 2368: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 2369: 	addi	%sp, %sp, 7
"01011000000000000010101000100100",	-- 2370: 	jal	yj_create_float_array
"10101011110111100000000000000111",	-- 2371: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 2372: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 2373: 	lli	%r2, 0
"00111100010111100000000000000110",	-- 2374: 	sw	%r2, [%sp + 6]
"00111100001111100000000000000111",	-- 2375: 	sw	%r1, [%sp + 7]
"00111111111111100000000000001000",	-- 2376: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 2377: 	addi	%sp, %sp, 9
"01011000000000000010101001000001",	-- 2378: 	jal	yj_read_float
"10101011110111100000000000001001",	-- 2379: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 2380: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000110",	-- 2381: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000111",	-- 2382: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 2383: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2384: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2385: 	lli	%r1, 1
"00111100001111100000000000001000",	-- 2386: 	sw	%r1, [%sp + 8]
"00111111111111100000000000001001",	-- 2387: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 2388: 	addi	%sp, %sp, 10
"01011000000000000010101001000001",	-- 2389: 	jal	yj_read_float
"10101011110111100000000000001010",	-- 2390: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 2391: 	lw	%ra, [%sp + 9]
"00111011110000010000000000001000",	-- 2392: 	lw	%r1, [%sp + 8]
"00111011110000100000000000000111",	-- 2393: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 2394: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2395: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2396: 	lli	%r1, 2
"00111100001111100000000000001001",	-- 2397: 	sw	%r1, [%sp + 9]
"00111111111111100000000000001010",	-- 2398: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 2399: 	addi	%sp, %sp, 11
"01011000000000000010101001000001",	-- 2400: 	jal	yj_read_float
"10101011110111100000000000001011",	-- 2401: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 2402: 	lw	%ra, [%sp + 10]
"00111011110000010000000000001001",	-- 2403: 	lw	%r1, [%sp + 9]
"00111011110000100000000000000111",	-- 2404: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 2405: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2406: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 2407: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 2408: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2409: 	lhif	%f0, 0.000000
"00111111111111100000000000001010",	-- 2410: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 2411: 	addi	%sp, %sp, 11
"01011000000000000010101000100100",	-- 2412: 	jal	yj_create_float_array
"10101011110111100000000000001011",	-- 2413: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 2414: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 2415: 	lli	%r2, 0
"00111100010111100000000000001010",	-- 2416: 	sw	%r2, [%sp + 10]
"00111100001111100000000000001011",	-- 2417: 	sw	%r1, [%sp + 11]
"00111111111111100000000000001100",	-- 2418: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 2419: 	addi	%sp, %sp, 13
"01011000000000000010101001000001",	-- 2420: 	jal	yj_read_float
"10101011110111100000000000001101",	-- 2421: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 2422: 	lw	%ra, [%sp + 12]
"00111011110000010000000000001010",	-- 2423: 	lw	%r1, [%sp + 10]
"00111011110000100000000000001011",	-- 2424: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 2425: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2426: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2427: 	lli	%r1, 1
"00111100001111100000000000001100",	-- 2428: 	sw	%r1, [%sp + 12]
"00111111111111100000000000001101",	-- 2429: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 2430: 	addi	%sp, %sp, 14
"01011000000000000010101001000001",	-- 2431: 	jal	yj_read_float
"10101011110111100000000000001110",	-- 2432: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 2433: 	lw	%ra, [%sp + 13]
"00111011110000010000000000001100",	-- 2434: 	lw	%r1, [%sp + 12]
"00111011110000100000000000001011",	-- 2435: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 2436: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2437: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2438: 	lli	%r1, 2
"00111100001111100000000000001101",	-- 2439: 	sw	%r1, [%sp + 13]
"00111111111111100000000000001110",	-- 2440: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 2441: 	addi	%sp, %sp, 15
"01011000000000000010101001000001",	-- 2442: 	jal	yj_read_float
"10101011110111100000000000001111",	-- 2443: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 2444: 	lw	%ra, [%sp + 14]
"00111011110000010000000000001101",	-- 2445: 	lw	%r1, [%sp + 13]
"00111011110000100000000000001011",	-- 2446: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 2447: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2448: 	sf	%f0, [%r1 + 0]
"00111111111111100000000000001110",	-- 2449: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 2450: 	addi	%sp, %sp, 15
"01011000000000000010101001000001",	-- 2451: 	jal	yj_read_float
"10101011110111100000000000001111",	-- 2452: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 2453: 	lw	%ra, [%sp + 14]
"00111111111111100000000000001110",	-- 2454: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 2455: 	addi	%sp, %sp, 15
"01011000000000000000010011011101",	-- 2456: 	jal	fisneg.2524
"10101011110111100000000000001111",	-- 2457: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 2458: 	lw	%ra, [%sp + 14]
"11001100000000100000000000000010",	-- 2459: 	lli	%r2, 2
"00010100000000000000000000000000",	-- 2460: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2461: 	lhif	%f0, 0.000000
"00111100001111100000000000001110",	-- 2462: 	sw	%r1, [%sp + 14]
"10000100000000100000100000000000",	-- 2463: 	add	%r1, %r0, %r2
"00111111111111100000000000001111",	-- 2464: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 2465: 	addi	%sp, %sp, 16
"01011000000000000010101000100100",	-- 2466: 	jal	yj_create_float_array
"10101011110111100000000000010000",	-- 2467: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 2468: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 2469: 	lli	%r2, 0
"00111100010111100000000000001111",	-- 2470: 	sw	%r2, [%sp + 15]
"00111100001111100000000000010000",	-- 2471: 	sw	%r1, [%sp + 16]
"00111111111111100000000000010001",	-- 2472: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 2473: 	addi	%sp, %sp, 18
"01011000000000000010101001000001",	-- 2474: 	jal	yj_read_float
"10101011110111100000000000010010",	-- 2475: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 2476: 	lw	%ra, [%sp + 17]
"00111011110000010000000000001111",	-- 2477: 	lw	%r1, [%sp + 15]
"00111011110000100000000000010000",	-- 2478: 	lw	%r2, [%sp + 16]
"10000100010000010000100000000000",	-- 2479: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2480: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2481: 	lli	%r1, 1
"00111100001111100000000000010001",	-- 2482: 	sw	%r1, [%sp + 17]
"00111111111111100000000000010010",	-- 2483: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 2484: 	addi	%sp, %sp, 19
"01011000000000000010101001000001",	-- 2485: 	jal	yj_read_float
"10101011110111100000000000010011",	-- 2486: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 2487: 	lw	%ra, [%sp + 18]
"00111011110000010000000000010001",	-- 2488: 	lw	%r1, [%sp + 17]
"00111011110000100000000000010000",	-- 2489: 	lw	%r2, [%sp + 16]
"10000100010000010000100000000000",	-- 2490: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2491: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 2492: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 2493: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2494: 	lhif	%f0, 0.000000
"00111111111111100000000000010010",	-- 2495: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 2496: 	addi	%sp, %sp, 19
"01011000000000000010101000100100",	-- 2497: 	jal	yj_create_float_array
"10101011110111100000000000010011",	-- 2498: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 2499: 	lw	%ra, [%sp + 18]
"11001100000000100000000000000000",	-- 2500: 	lli	%r2, 0
"00111100010111100000000000010010",	-- 2501: 	sw	%r2, [%sp + 18]
"00111100001111100000000000010011",	-- 2502: 	sw	%r1, [%sp + 19]
"00111111111111100000000000010100",	-- 2503: 	sw	%ra, [%sp + 20]
"10100111110111100000000000010101",	-- 2504: 	addi	%sp, %sp, 21
"01011000000000000010101001000001",	-- 2505: 	jal	yj_read_float
"10101011110111100000000000010101",	-- 2506: 	subi	%sp, %sp, 21
"00111011110111110000000000010100",	-- 2507: 	lw	%ra, [%sp + 20]
"00111011110000010000000000010010",	-- 2508: 	lw	%r1, [%sp + 18]
"00111011110000100000000000010011",	-- 2509: 	lw	%r2, [%sp + 19]
"10000100010000010000100000000000",	-- 2510: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2511: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2512: 	lli	%r1, 1
"00111100001111100000000000010100",	-- 2513: 	sw	%r1, [%sp + 20]
"00111111111111100000000000010101",	-- 2514: 	sw	%ra, [%sp + 21]
"10100111110111100000000000010110",	-- 2515: 	addi	%sp, %sp, 22
"01011000000000000010101001000001",	-- 2516: 	jal	yj_read_float
"10101011110111100000000000010110",	-- 2517: 	subi	%sp, %sp, 22
"00111011110111110000000000010101",	-- 2518: 	lw	%ra, [%sp + 21]
"00111011110000010000000000010100",	-- 2519: 	lw	%r1, [%sp + 20]
"00111011110000100000000000010011",	-- 2520: 	lw	%r2, [%sp + 19]
"10000100010000010000100000000000",	-- 2521: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2522: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2523: 	lli	%r1, 2
"00111100001111100000000000010101",	-- 2524: 	sw	%r1, [%sp + 21]
"00111111111111100000000000010110",	-- 2525: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 2526: 	addi	%sp, %sp, 23
"01011000000000000010101001000001",	-- 2527: 	jal	yj_read_float
"10101011110111100000000000010111",	-- 2528: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 2529: 	lw	%ra, [%sp + 22]
"00111011110000010000000000010101",	-- 2530: 	lw	%r1, [%sp + 21]
"00111011110000100000000000010011",	-- 2531: 	lw	%r2, [%sp + 19]
"10000100010000010000100000000000",	-- 2532: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2533: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 2534: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 2535: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2536: 	lhif	%f0, 0.000000
"00111111111111100000000000010110",	-- 2537: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 2538: 	addi	%sp, %sp, 23
"01011000000000000010101000100100",	-- 2539: 	jal	yj_create_float_array
"10101011110111100000000000010111",	-- 2540: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 2541: 	lw	%ra, [%sp + 22]
"11001100000000100000000000000000",	-- 2542: 	lli	%r2, 0
"00111011110000110000000000000101",	-- 2543: 	lw	%r3, [%sp + 5]
"00111100001111100000000000010110",	-- 2544: 	sw	%r1, [%sp + 22]
"00101000011000100000000000000010",	-- 2545: 	bneq	%r3, %r2, bneq_else.8962
"01010100000000000000101000100011",	-- 2546: 	j	bneq_cont.8963
	-- bneq_else.8962:
"11001100000000100000000000000000",	-- 2547: 	lli	%r2, 0
"00111100010111100000000000010111",	-- 2548: 	sw	%r2, [%sp + 23]
"00111111111111100000000000011000",	-- 2549: 	sw	%ra, [%sp + 24]
"10100111110111100000000000011001",	-- 2550: 	addi	%sp, %sp, 25
"01011000000000000010101001000001",	-- 2551: 	jal	yj_read_float
"10101011110111100000000000011001",	-- 2552: 	subi	%sp, %sp, 25
"00111011110111110000000000011000",	-- 2553: 	lw	%ra, [%sp + 24]
"00111111111111100000000000011000",	-- 2554: 	sw	%ra, [%sp + 24]
"10100111110111100000000000011001",	-- 2555: 	addi	%sp, %sp, 25
"01011000000000000000011011000110",	-- 2556: 	jal	rad.2693
"10101011110111100000000000011001",	-- 2557: 	subi	%sp, %sp, 25
"00111011110111110000000000011000",	-- 2558: 	lw	%ra, [%sp + 24]
"00111011110000010000000000010111",	-- 2559: 	lw	%r1, [%sp + 23]
"00111011110000100000000000010110",	-- 2560: 	lw	%r2, [%sp + 22]
"10000100010000010000100000000000",	-- 2561: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2562: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2563: 	lli	%r1, 1
"00111100001111100000000000011000",	-- 2564: 	sw	%r1, [%sp + 24]
"00111111111111100000000000011001",	-- 2565: 	sw	%ra, [%sp + 25]
"10100111110111100000000000011010",	-- 2566: 	addi	%sp, %sp, 26
"01011000000000000010101001000001",	-- 2567: 	jal	yj_read_float
"10101011110111100000000000011010",	-- 2568: 	subi	%sp, %sp, 26
"00111011110111110000000000011001",	-- 2569: 	lw	%ra, [%sp + 25]
"00111111111111100000000000011001",	-- 2570: 	sw	%ra, [%sp + 25]
"10100111110111100000000000011010",	-- 2571: 	addi	%sp, %sp, 26
"01011000000000000000011011000110",	-- 2572: 	jal	rad.2693
"10101011110111100000000000011010",	-- 2573: 	subi	%sp, %sp, 26
"00111011110111110000000000011001",	-- 2574: 	lw	%ra, [%sp + 25]
"00111011110000010000000000011000",	-- 2575: 	lw	%r1, [%sp + 24]
"00111011110000100000000000010110",	-- 2576: 	lw	%r2, [%sp + 22]
"10000100010000010000100000000000",	-- 2577: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2578: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2579: 	lli	%r1, 2
"00111100001111100000000000011001",	-- 2580: 	sw	%r1, [%sp + 25]
"00111111111111100000000000011010",	-- 2581: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 2582: 	addi	%sp, %sp, 27
"01011000000000000010101001000001",	-- 2583: 	jal	yj_read_float
"10101011110111100000000000011011",	-- 2584: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 2585: 	lw	%ra, [%sp + 26]
"00111111111111100000000000011010",	-- 2586: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 2587: 	addi	%sp, %sp, 27
"01011000000000000000011011000110",	-- 2588: 	jal	rad.2693
"10101011110111100000000000011011",	-- 2589: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 2590: 	lw	%ra, [%sp + 26]
"00111011110000010000000000011001",	-- 2591: 	lw	%r1, [%sp + 25]
"00111011110000100000000000010110",	-- 2592: 	lw	%r2, [%sp + 22]
"10000100010000010000100000000000",	-- 2593: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2594: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.8963:
"11001100000000010000000000000010",	-- 2595: 	lli	%r1, 2
"00111011110000100000000000000011",	-- 2596: 	lw	%r2, [%sp + 3]
"00101000010000010000000000000011",	-- 2597: 	bneq	%r2, %r1, bneq_else.8964
"11001100000000010000000000000001",	-- 2598: 	lli	%r1, 1
"01010100000000000000101000101001",	-- 2599: 	j	bneq_cont.8965
	-- bneq_else.8964:
"00111011110000010000000000001110",	-- 2600: 	lw	%r1, [%sp + 14]
	-- bneq_cont.8965:
"11001100000000110000000000000100",	-- 2601: 	lli	%r3, 4
"00010100000000000000000000000000",	-- 2602: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2603: 	lhif	%f0, 0.000000
"00111100001111100000000000011010",	-- 2604: 	sw	%r1, [%sp + 26]
"10000100000000110000100000000000",	-- 2605: 	add	%r1, %r0, %r3
"00111111111111100000000000011011",	-- 2606: 	sw	%ra, [%sp + 27]
"10100111110111100000000000011100",	-- 2607: 	addi	%sp, %sp, 28
"01011000000000000010101000100100",	-- 2608: 	jal	yj_create_float_array
"10101011110111100000000000011100",	-- 2609: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 2610: 	lw	%ra, [%sp + 27]
"10000100000111010001000000000000",	-- 2611: 	add	%r2, %r0, %hp
"10100111101111010000000000001011",	-- 2612: 	addi	%hp, %hp, 11
"00111100001000100000000000001010",	-- 2613: 	sw	%r1, [%r2 + 10]
"00111011110000010000000000010110",	-- 2614: 	lw	%r1, [%sp + 22]
"00111100001000100000000000001001",	-- 2615: 	sw	%r1, [%r2 + 9]
"00111011110000110000000000010011",	-- 2616: 	lw	%r3, [%sp + 19]
"00111100011000100000000000001000",	-- 2617: 	sw	%r3, [%r2 + 8]
"00111011110000110000000000010000",	-- 2618: 	lw	%r3, [%sp + 16]
"00111100011000100000000000000111",	-- 2619: 	sw	%r3, [%r2 + 7]
"00111011110000110000000000011010",	-- 2620: 	lw	%r3, [%sp + 26]
"00111100011000100000000000000110",	-- 2621: 	sw	%r3, [%r2 + 6]
"00111011110000110000000000001011",	-- 2622: 	lw	%r3, [%sp + 11]
"00111100011000100000000000000101",	-- 2623: 	sw	%r3, [%r2 + 5]
"00111011110000110000000000000111",	-- 2624: 	lw	%r3, [%sp + 7]
"00111100011000100000000000000100",	-- 2625: 	sw	%r3, [%r2 + 4]
"00111011110001000000000000000101",	-- 2626: 	lw	%r4, [%sp + 5]
"00111100100000100000000000000011",	-- 2627: 	sw	%r4, [%r2 + 3]
"00111011110001010000000000000100",	-- 2628: 	lw	%r5, [%sp + 4]
"00111100101000100000000000000010",	-- 2629: 	sw	%r5, [%r2 + 2]
"00111011110001010000000000000011",	-- 2630: 	lw	%r5, [%sp + 3]
"00111100101000100000000000000001",	-- 2631: 	sw	%r5, [%r2 + 1]
"00111011110001100000000000000010",	-- 2632: 	lw	%r6, [%sp + 2]
"00111100110000100000000000000000",	-- 2633: 	sw	%r6, [%r2 + 0]
"00111011110001100000000000000000",	-- 2634: 	lw	%r6, [%sp + 0]
"00111011110001110000000000000001",	-- 2635: 	lw	%r7, [%sp + 1]
"10000100111001100011000000000000",	-- 2636: 	add	%r6, %r7, %r6
"00111100010001100000000000000000",	-- 2637: 	sw	%r2, [%r6 + 0]
"11001100000000100000000000000011",	-- 2638: 	lli	%r2, 3
"00101000101000100000000001101110",	-- 2639: 	bneq	%r5, %r2, bneq_else.8966
"11001100000000100000000000000000",	-- 2640: 	lli	%r2, 0
"10000100011000100001000000000000",	-- 2641: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 2642: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000000",	-- 2643: 	lli	%r2, 0
"00111100010111100000000000011011",	-- 2644: 	sw	%r2, [%sp + 27]
"10110000000111100000000000011100",	-- 2645: 	sf	%f0, [%sp + 28]
"00111111111111100000000000011101",	-- 2646: 	sw	%ra, [%sp + 29]
"10100111110111100000000000011110",	-- 2647: 	addi	%sp, %sp, 30
"01011000000000000000010011100100",	-- 2648: 	jal	fiszero.2526
"10101011110111100000000000011110",	-- 2649: 	subi	%sp, %sp, 30
"00111011110111110000000000011101",	-- 2650: 	lw	%ra, [%sp + 29]
"11001100000000100000000000000000",	-- 2651: 	lli	%r2, 0
"00101000001000100000000000010010",	-- 2652: 	bneq	%r1, %r2, bneq_else.8968
"10010011110000000000000000011100",	-- 2653: 	lf	%f0, [%sp + 28]
"00111111111111100000000000011101",	-- 2654: 	sw	%ra, [%sp + 29]
"10100111110111100000000000011110",	-- 2655: 	addi	%sp, %sp, 30
"01011000000000000000010100000010",	-- 2656: 	jal	sgn.2568
"10101011110111100000000000011110",	-- 2657: 	subi	%sp, %sp, 30
"00111011110111110000000000011101",	-- 2658: 	lw	%ra, [%sp + 29]
"10010011110000010000000000011100",	-- 2659: 	lf	%f1, [%sp + 28]
"10110000000111100000000000011101",	-- 2660: 	sf	%f0, [%sp + 29]
"00001100001000000000000000000000",	-- 2661: 	movf	%f0, %f1
"00111111111111100000000000011110",	-- 2662: 	sw	%ra, [%sp + 30]
"10100111110111100000000000011111",	-- 2663: 	addi	%sp, %sp, 31
"01011000000000000000010011110001",	-- 2664: 	jal	fsqr.2530
"10101011110111100000000000011111",	-- 2665: 	subi	%sp, %sp, 31
"00111011110111110000000000011110",	-- 2666: 	lw	%ra, [%sp + 30]
"10010011110000010000000000011101",	-- 2667: 	lf	%f1, [%sp + 29]
"11101100001000000000000000000000",	-- 2668: 	divf	%f0, %f1, %f0
"01010100000000000000101001110000",	-- 2669: 	j	bneq_cont.8969
	-- bneq_else.8968:
"00010100000000000000000000000000",	-- 2670: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2671: 	lhif	%f0, 0.000000
	-- bneq_cont.8969:
"00111011110000010000000000011011",	-- 2672: 	lw	%r1, [%sp + 27]
"00111011110000100000000000000111",	-- 2673: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 2674: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2675: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2676: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 2677: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 2678: 	lf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 2679: 	lli	%r1, 1
"00111100001111100000000000011110",	-- 2680: 	sw	%r1, [%sp + 30]
"10110000000111100000000000011111",	-- 2681: 	sf	%f0, [%sp + 31]
"00111111111111100000000000100000",	-- 2682: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 2683: 	addi	%sp, %sp, 33
"01011000000000000000010011100100",	-- 2684: 	jal	fiszero.2526
"10101011110111100000000000100001",	-- 2685: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 2686: 	lw	%ra, [%sp + 32]
"11001100000000100000000000000000",	-- 2687: 	lli	%r2, 0
"00101000001000100000000000010010",	-- 2688: 	bneq	%r1, %r2, bneq_else.8970
"10010011110000000000000000011111",	-- 2689: 	lf	%f0, [%sp + 31]
"00111111111111100000000000100000",	-- 2690: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 2691: 	addi	%sp, %sp, 33
"01011000000000000000010100000010",	-- 2692: 	jal	sgn.2568
"10101011110111100000000000100001",	-- 2693: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 2694: 	lw	%ra, [%sp + 32]
"10010011110000010000000000011111",	-- 2695: 	lf	%f1, [%sp + 31]
"10110000000111100000000000100000",	-- 2696: 	sf	%f0, [%sp + 32]
"00001100001000000000000000000000",	-- 2697: 	movf	%f0, %f1
"00111111111111100000000000100001",	-- 2698: 	sw	%ra, [%sp + 33]
"10100111110111100000000000100010",	-- 2699: 	addi	%sp, %sp, 34
"01011000000000000000010011110001",	-- 2700: 	jal	fsqr.2530
"10101011110111100000000000100010",	-- 2701: 	subi	%sp, %sp, 34
"00111011110111110000000000100001",	-- 2702: 	lw	%ra, [%sp + 33]
"10010011110000010000000000100000",	-- 2703: 	lf	%f1, [%sp + 32]
"11101100001000000000000000000000",	-- 2704: 	divf	%f0, %f1, %f0
"01010100000000000000101010010100",	-- 2705: 	j	bneq_cont.8971
	-- bneq_else.8970:
"00010100000000000000000000000000",	-- 2706: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2707: 	lhif	%f0, 0.000000
	-- bneq_cont.8971:
"00111011110000010000000000011110",	-- 2708: 	lw	%r1, [%sp + 30]
"00111011110000100000000000000111",	-- 2709: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 2710: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2711: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2712: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 2713: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 2714: 	lf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 2715: 	lli	%r1, 2
"00111100001111100000000000100001",	-- 2716: 	sw	%r1, [%sp + 33]
"10110000000111100000000000100010",	-- 2717: 	sf	%f0, [%sp + 34]
"00111111111111100000000000100011",	-- 2718: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 2719: 	addi	%sp, %sp, 36
"01011000000000000000010011100100",	-- 2720: 	jal	fiszero.2526
"10101011110111100000000000100100",	-- 2721: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 2722: 	lw	%ra, [%sp + 35]
"11001100000000100000000000000000",	-- 2723: 	lli	%r2, 0
"00101000001000100000000000010010",	-- 2724: 	bneq	%r1, %r2, bneq_else.8972
"10010011110000000000000000100010",	-- 2725: 	lf	%f0, [%sp + 34]
"00111111111111100000000000100011",	-- 2726: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 2727: 	addi	%sp, %sp, 36
"01011000000000000000010100000010",	-- 2728: 	jal	sgn.2568
"10101011110111100000000000100100",	-- 2729: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 2730: 	lw	%ra, [%sp + 35]
"10010011110000010000000000100010",	-- 2731: 	lf	%f1, [%sp + 34]
"10110000000111100000000000100011",	-- 2732: 	sf	%f0, [%sp + 35]
"00001100001000000000000000000000",	-- 2733: 	movf	%f0, %f1
"00111111111111100000000000100100",	-- 2734: 	sw	%ra, [%sp + 36]
"10100111110111100000000000100101",	-- 2735: 	addi	%sp, %sp, 37
"01011000000000000000010011110001",	-- 2736: 	jal	fsqr.2530
"10101011110111100000000000100101",	-- 2737: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 2738: 	lw	%ra, [%sp + 36]
"10010011110000010000000000100011",	-- 2739: 	lf	%f1, [%sp + 35]
"11101100001000000000000000000000",	-- 2740: 	divf	%f0, %f1, %f0
"01010100000000000000101010111000",	-- 2741: 	j	bneq_cont.8973
	-- bneq_else.8972:
"00010100000000000000000000000000",	-- 2742: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 2743: 	lhif	%f0, 0.000000
	-- bneq_cont.8973:
"00111011110000010000000000100001",	-- 2744: 	lw	%r1, [%sp + 33]
"00111011110000100000000000000111",	-- 2745: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 2746: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 2747: 	sf	%f0, [%r1 + 0]
"01010100000000000000101011001100",	-- 2748: 	j	bneq_cont.8967
	-- bneq_else.8966:
"11001100000000100000000000000010",	-- 2749: 	lli	%r2, 2
"00101000101000100000000000001110",	-- 2750: 	bneq	%r5, %r2, bneq_else.8974
"11001100000000100000000000000000",	-- 2751: 	lli	%r2, 0
"00111011110001010000000000001110",	-- 2752: 	lw	%r5, [%sp + 14]
"00101000101000100000000000000011",	-- 2753: 	bneq	%r5, %r2, bneq_else.8976
"11001100000000100000000000000001",	-- 2754: 	lli	%r2, 1
"01010100000000000000101011000101",	-- 2755: 	j	bneq_cont.8977
	-- bneq_else.8976:
"11001100000000100000000000000000",	-- 2756: 	lli	%r2, 0
	-- bneq_cont.8977:
"10000100000000110000100000000000",	-- 2757: 	add	%r1, %r0, %r3
"00111111111111100000000000100100",	-- 2758: 	sw	%ra, [%sp + 36]
"10100111110111100000000000100101",	-- 2759: 	addi	%sp, %sp, 37
"01011000000000000000010101010000",	-- 2760: 	jal	vecunit_sgn.2594
"10101011110111100000000000100101",	-- 2761: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 2762: 	lw	%ra, [%sp + 36]
"01010100000000000000101011001100",	-- 2763: 	j	bneq_cont.8975
	-- bneq_else.8974:
	-- bneq_cont.8975:
	-- bneq_cont.8967:
"11001100000000010000000000000000",	-- 2764: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 2765: 	lw	%r2, [%sp + 5]
"00101000010000010000000000000010",	-- 2766: 	bneq	%r2, %r1, bneq_else.8978
"01010100000000000000101011010111",	-- 2767: 	j	bneq_cont.8979
	-- bneq_else.8978:
"00111011110000010000000000000111",	-- 2768: 	lw	%r1, [%sp + 7]
"00111011110000100000000000010110",	-- 2769: 	lw	%r2, [%sp + 22]
"00111111111111100000000000100100",	-- 2770: 	sw	%ra, [%sp + 36]
"10100111110111100000000000100101",	-- 2771: 	addi	%sp, %sp, 37
"01011000000000000000011111111001",	-- 2772: 	jal	rotate_quadratic_matrix.2699
"10101011110111100000000000100101",	-- 2773: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 2774: 	lw	%ra, [%sp + 36]
	-- bneq_cont.8979:
"11001100000000010000000000000001",	-- 2775: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 2776: 	jr	%ra
	-- read_object.2704:
"00111011011000100000000000000010",	-- 2777: 	lw	%r2, [%r27 + 2]
"00111011011000110000000000000001",	-- 2778: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000111100",	-- 2779: 	lli	%r4, 60
"00110000100000010000000000000010",	-- 2780: 	bgt	%r4, %r1, bgt_else.8980
"01001111111000000000000000000000",	-- 2781: 	jr	%ra
	-- bgt_else.8980:
"00111111011111100000000000000000",	-- 2782: 	sw	%r27, [%sp + 0]
"00111100001111100000000000000001",	-- 2783: 	sw	%r1, [%sp + 1]
"00111100011111100000000000000010",	-- 2784: 	sw	%r3, [%sp + 2]
"10000100000000101101100000000000",	-- 2785: 	add	%r27, %r0, %r2
"00111111111111100000000000000011",	-- 2786: 	sw	%ra, [%sp + 3]
"00111011011110100000000000000000",	-- 2787: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000100",	-- 2788: 	addi	%sp, %sp, 4
"01010011010000000000000000000000",	-- 2789: 	jalr	%r26
"10101011110111100000000000000100",	-- 2790: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 2791: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000000",	-- 2792: 	lli	%r2, 0
"00101000001000100000000000000111",	-- 2793: 	bneq	%r1, %r2, bneq_else.8982
"11001100000000010000000000000000",	-- 2794: 	lli	%r1, 0
"00111011110000100000000000000010",	-- 2795: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 2796: 	add	%r1, %r2, %r1
"00111011110000100000000000000001",	-- 2797: 	lw	%r2, [%sp + 1]
"00111100010000010000000000000000",	-- 2798: 	sw	%r2, [%r1 + 0]
"01001111111000000000000000000000",	-- 2799: 	jr	%ra
	-- bneq_else.8982:
"11001100000000010000000000000001",	-- 2800: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 2801: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 2802: 	add	%r1, %r2, %r1
"00111011110110110000000000000000",	-- 2803: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 2804: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 2805: 	jr	%r26
	-- read_all_object.2706:
"00111011011110110000000000000001",	-- 2806: 	lw	%r27, [%r27 + 1]
"11001100000000010000000000000000",	-- 2807: 	lli	%r1, 0
"00111011011110100000000000000000",	-- 2808: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 2809: 	jr	%r26
	-- read_net_item.2708:
"00111100001111100000000000000000",	-- 2810: 	sw	%r1, [%sp + 0]
"00111111111111100000000000000001",	-- 2811: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 2812: 	addi	%sp, %sp, 2
"01011000000000000010101000110100",	-- 2813: 	jal	yj_read_int
"10101011110111100000000000000010",	-- 2814: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 2815: 	lw	%ra, [%sp + 1]
"11001100000000101111111111111111",	-- 2816: 	lli	%r2, -1
"11001000000000101111111111111111",	-- 2817: 	lhi	%r2, -1
"00101000001000100000000000000111",	-- 2818: 	bneq	%r1, %r2, bneq_else.8984
"11001100000000010000000000000001",	-- 2819: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 2820: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 2821: 	add	%r1, %r2, %r1
"11001100000000101111111111111111",	-- 2822: 	lli	%r2, -1
"11001000000000101111111111111111",	-- 2823: 	lhi	%r2, -1
"01010100000000000010101000011100",	-- 2824: 	j	yj_create_array
	-- bneq_else.8984:
"11001100000000100000000000000001",	-- 2825: 	lli	%r2, 1
"00111011110000110000000000000000",	-- 2826: 	lw	%r3, [%sp + 0]
"10000100011000100001000000000000",	-- 2827: 	add	%r2, %r3, %r2
"00111100001111100000000000000001",	-- 2828: 	sw	%r1, [%sp + 1]
"10000100000000100000100000000000",	-- 2829: 	add	%r1, %r0, %r2
"00111111111111100000000000000010",	-- 2830: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 2831: 	addi	%sp, %sp, 3
"01011000000000000000101011111010",	-- 2832: 	jal	read_net_item.2708
"10101011110111100000000000000011",	-- 2833: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 2834: 	lw	%ra, [%sp + 2]
"00111011110000100000000000000000",	-- 2835: 	lw	%r2, [%sp + 0]
"10000100001000100001000000000000",	-- 2836: 	add	%r2, %r1, %r2
"00111011110000110000000000000001",	-- 2837: 	lw	%r3, [%sp + 1]
"00111100011000100000000000000000",	-- 2838: 	sw	%r3, [%r2 + 0]
"01001111111000000000000000000000",	-- 2839: 	jr	%ra
	-- read_or_network.2710:
"11001100000000100000000000000000",	-- 2840: 	lli	%r2, 0
"00111100001111100000000000000000",	-- 2841: 	sw	%r1, [%sp + 0]
"10000100000000100000100000000000",	-- 2842: 	add	%r1, %r0, %r2
"00111111111111100000000000000001",	-- 2843: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 2844: 	addi	%sp, %sp, 2
"01011000000000000000101011111010",	-- 2845: 	jal	read_net_item.2708
"10101011110111100000000000000010",	-- 2846: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 2847: 	lw	%ra, [%sp + 1]
"10000100000000010001000000000000",	-- 2848: 	add	%r2, %r0, %r1
"11001100000000010000000000000000",	-- 2849: 	lli	%r1, 0
"10000100010000010000100000000000",	-- 2850: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 2851: 	lw	%r1, [%r1 + 0]
"11001100000000111111111111111111",	-- 2852: 	lli	%r3, -1
"11001000000000111111111111111111",	-- 2853: 	lhi	%r3, -1
"00101000001000110000000000000101",	-- 2854: 	bneq	%r1, %r3, bneq_else.8985
"11001100000000010000000000000001",	-- 2855: 	lli	%r1, 1
"00111011110000110000000000000000",	-- 2856: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 2857: 	add	%r1, %r3, %r1
"01010100000000000010101000011100",	-- 2858: 	j	yj_create_array
	-- bneq_else.8985:
"11001100000000010000000000000001",	-- 2859: 	lli	%r1, 1
"00111011110000110000000000000000",	-- 2860: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 2861: 	add	%r1, %r3, %r1
"00111100010111100000000000000001",	-- 2862: 	sw	%r2, [%sp + 1]
"00111111111111100000000000000010",	-- 2863: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 2864: 	addi	%sp, %sp, 3
"01011000000000000000101100011000",	-- 2865: 	jal	read_or_network.2710
"10101011110111100000000000000011",	-- 2866: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 2867: 	lw	%ra, [%sp + 2]
"00111011110000100000000000000000",	-- 2868: 	lw	%r2, [%sp + 0]
"10000100001000100001000000000000",	-- 2869: 	add	%r2, %r1, %r2
"00111011110000110000000000000001",	-- 2870: 	lw	%r3, [%sp + 1]
"00111100011000100000000000000000",	-- 2871: 	sw	%r3, [%r2 + 0]
"01001111111000000000000000000000",	-- 2872: 	jr	%ra
	-- read_and_network.2712:
"00111011011000100000000000000001",	-- 2873: 	lw	%r2, [%r27 + 1]
"11001100000000110000000000000000",	-- 2874: 	lli	%r3, 0
"00111111011111100000000000000000",	-- 2875: 	sw	%r27, [%sp + 0]
"00111100001111100000000000000001",	-- 2876: 	sw	%r1, [%sp + 1]
"00111100010111100000000000000010",	-- 2877: 	sw	%r2, [%sp + 2]
"10000100000000110000100000000000",	-- 2878: 	add	%r1, %r0, %r3
"00111111111111100000000000000011",	-- 2879: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 2880: 	addi	%sp, %sp, 4
"01011000000000000000101011111010",	-- 2881: 	jal	read_net_item.2708
"10101011110111100000000000000100",	-- 2882: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 2883: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000000",	-- 2884: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 2885: 	add	%r2, %r1, %r2
"00111000010000100000000000000000",	-- 2886: 	lw	%r2, [%r2 + 0]
"11001100000000111111111111111111",	-- 2887: 	lli	%r3, -1
"11001000000000111111111111111111",	-- 2888: 	lhi	%r3, -1
"00101000010000110000000000000010",	-- 2889: 	bneq	%r2, %r3, bneq_else.8986
"01001111111000000000000000000000",	-- 2890: 	jr	%ra
	-- bneq_else.8986:
"00111011110000100000000000000001",	-- 2891: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000010",	-- 2892: 	lw	%r3, [%sp + 2]
"10000100011000100001100000000000",	-- 2893: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 2894: 	sw	%r1, [%r3 + 0]
"11001100000000010000000000000001",	-- 2895: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 2896: 	add	%r1, %r2, %r1
"00111011110110110000000000000000",	-- 2897: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 2898: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 2899: 	jr	%r26
	-- read_parameter.2714:
"00111011011000010000000000000101",	-- 2900: 	lw	%r1, [%r27 + 5]
"00111011011000100000000000000100",	-- 2901: 	lw	%r2, [%r27 + 4]
"00111011011000110000000000000011",	-- 2902: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 2903: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 2904: 	lw	%r5, [%r27 + 1]
"00111100101111100000000000000000",	-- 2905: 	sw	%r5, [%sp + 0]
"00111100011111100000000000000001",	-- 2906: 	sw	%r3, [%sp + 1]
"00111100100111100000000000000010",	-- 2907: 	sw	%r4, [%sp + 2]
"00111100010111100000000000000011",	-- 2908: 	sw	%r2, [%sp + 3]
"10000100000000011101100000000000",	-- 2909: 	add	%r27, %r0, %r1
"00111111111111100000000000000100",	-- 2910: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 2911: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 2912: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 2913: 	jalr	%r26
"10101011110111100000000000000101",	-- 2914: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 2915: 	lw	%ra, [%sp + 4]
"00111011110110110000000000000011",	-- 2916: 	lw	%r27, [%sp + 3]
"00111111111111100000000000000100",	-- 2917: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 2918: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 2919: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 2920: 	jalr	%r26
"10101011110111100000000000000101",	-- 2921: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 2922: 	lw	%ra, [%sp + 4]
"00111011110110110000000000000010",	-- 2923: 	lw	%r27, [%sp + 2]
"00111111111111100000000000000100",	-- 2924: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 2925: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 2926: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 2927: 	jalr	%r26
"10101011110111100000000000000101",	-- 2928: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 2929: 	lw	%ra, [%sp + 4]
"11001100000000010000000000000000",	-- 2930: 	lli	%r1, 0
"00111011110110110000000000000001",	-- 2931: 	lw	%r27, [%sp + 1]
"00111111111111100000000000000100",	-- 2932: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 2933: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 2934: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 2935: 	jalr	%r26
"10101011110111100000000000000101",	-- 2936: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 2937: 	lw	%ra, [%sp + 4]
"11001100000000010000000000000000",	-- 2938: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 2939: 	lli	%r2, 0
"00111100001111100000000000000100",	-- 2940: 	sw	%r1, [%sp + 4]
"10000100000000100000100000000000",	-- 2941: 	add	%r1, %r0, %r2
"00111111111111100000000000000101",	-- 2942: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 2943: 	addi	%sp, %sp, 6
"01011000000000000000101100011000",	-- 2944: 	jal	read_or_network.2710
"10101011110111100000000000000110",	-- 2945: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 2946: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000100",	-- 2947: 	lw	%r2, [%sp + 4]
"00111011110000110000000000000000",	-- 2948: 	lw	%r3, [%sp + 0]
"10000100011000100001000000000000",	-- 2949: 	add	%r2, %r3, %r2
"00111100001000100000000000000000",	-- 2950: 	sw	%r1, [%r2 + 0]
"01001111111000000000000000000000",	-- 2951: 	jr	%ra
	-- solver_rect_surface.2716:
"00111011011001100000000000000001",	-- 2952: 	lw	%r6, [%r27 + 1]
"10000100010000110011100000000000",	-- 2953: 	add	%r7, %r2, %r3
"10010000111000110000000000000000",	-- 2954: 	lf	%f3, [%r7 + 0]
"00111100110111100000000000000000",	-- 2955: 	sw	%r6, [%sp + 0]
"10110000010111100000000000000001",	-- 2956: 	sf	%f2, [%sp + 1]
"00111100101111100000000000000010",	-- 2957: 	sw	%r5, [%sp + 2]
"10110000001111100000000000000011",	-- 2958: 	sf	%f1, [%sp + 3]
"00111100100111100000000000000100",	-- 2959: 	sw	%r4, [%sp + 4]
"10110000000111100000000000000101",	-- 2960: 	sf	%f0, [%sp + 5]
"00111100011111100000000000000110",	-- 2961: 	sw	%r3, [%sp + 6]
"00111100010111100000000000000111",	-- 2962: 	sw	%r2, [%sp + 7]
"00111100001111100000000000001000",	-- 2963: 	sw	%r1, [%sp + 8]
"00001100011000000000000000000000",	-- 2964: 	movf	%f0, %f3
"00111111111111100000000000001001",	-- 2965: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 2966: 	addi	%sp, %sp, 10
"01011000000000000000010011100100",	-- 2967: 	jal	fiszero.2526
"10101011110111100000000000001010",	-- 2968: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 2969: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000000",	-- 2970: 	lli	%r2, 0
"00101000001000100000000001101011",	-- 2971: 	bneq	%r1, %r2, bneq_else.8989
"00111011110000010000000000001000",	-- 2972: 	lw	%r1, [%sp + 8]
"00111111111111100000000000001001",	-- 2973: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 2974: 	addi	%sp, %sp, 10
"01011000000000000000011001101001",	-- 2975: 	jal	o_param_abc.2638
"10101011110111100000000000001010",	-- 2976: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 2977: 	lw	%ra, [%sp + 9]
"00111011110000100000000000001000",	-- 2978: 	lw	%r2, [%sp + 8]
"00111100001111100000000000001001",	-- 2979: 	sw	%r1, [%sp + 9]
"10000100000000100000100000000000",	-- 2980: 	add	%r1, %r0, %r2
"00111111111111100000000000001010",	-- 2981: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 2982: 	addi	%sp, %sp, 11
"01011000000000000000011001010110",	-- 2983: 	jal	o_isinvert.2628
"10101011110111100000000000001011",	-- 2984: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 2985: 	lw	%ra, [%sp + 10]
"00111011110000100000000000000110",	-- 2986: 	lw	%r2, [%sp + 6]
"00111011110000110000000000000111",	-- 2987: 	lw	%r3, [%sp + 7]
"10000100011000100010000000000000",	-- 2988: 	add	%r4, %r3, %r2
"10010000100000000000000000000000",	-- 2989: 	lf	%f0, [%r4 + 0]
"00111100001111100000000000001010",	-- 2990: 	sw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 2991: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 2992: 	addi	%sp, %sp, 12
"01011000000000000000010011011101",	-- 2993: 	jal	fisneg.2524
"10101011110111100000000000001100",	-- 2994: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 2995: 	lw	%ra, [%sp + 11]
"10000100000000010001000000000000",	-- 2996: 	add	%r2, %r0, %r1
"00111011110000010000000000001010",	-- 2997: 	lw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 2998: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 2999: 	addi	%sp, %sp, 12
"01011000000000000000010011111000",	-- 3000: 	jal	xor.2565
"10101011110111100000000000001100",	-- 3001: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3002: 	lw	%ra, [%sp + 11]
"00111011110000100000000000000110",	-- 3003: 	lw	%r2, [%sp + 6]
"00111011110000110000000000001001",	-- 3004: 	lw	%r3, [%sp + 9]
"10000100011000100010000000000000",	-- 3005: 	add	%r4, %r3, %r2
"10010000100000000000000000000000",	-- 3006: 	lf	%f0, [%r4 + 0]
"00111111111111100000000000001011",	-- 3007: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 3008: 	addi	%sp, %sp, 12
"01011000000000000000010100011011",	-- 3009: 	jal	fneg_cond.2570
"10101011110111100000000000001100",	-- 3010: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3011: 	lw	%ra, [%sp + 11]
"10010011110000010000000000000101",	-- 3012: 	lf	%f1, [%sp + 5]
"11100100000000010000000000000000",	-- 3013: 	subf	%f0, %f0, %f1
"00111011110000010000000000000110",	-- 3014: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000111",	-- 3015: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 3016: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3017: 	lf	%f1, [%r1 + 0]
"11101100000000010000000000000000",	-- 3018: 	divf	%f0, %f0, %f1
"00111011110000010000000000000100",	-- 3019: 	lw	%r1, [%sp + 4]
"10000100010000010001100000000000",	-- 3020: 	add	%r3, %r2, %r1
"10010000011000010000000000000000",	-- 3021: 	lf	%f1, [%r3 + 0]
"11101000000000010000100000000000",	-- 3022: 	mulf	%f1, %f0, %f1
"10010011110000100000000000000011",	-- 3023: 	lf	%f2, [%sp + 3]
"11100000001000100000100000000000",	-- 3024: 	addf	%f1, %f1, %f2
"10110000000111100000000000001011",	-- 3025: 	sf	%f0, [%sp + 11]
"00001100001000000000000000000000",	-- 3026: 	movf	%f0, %f1
"00111111111111100000000000001100",	-- 3027: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3028: 	addi	%sp, %sp, 13
"01011000000000000010101001001111",	-- 3029: 	jal	yj_fabs
"10101011110111100000000000001101",	-- 3030: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3031: 	lw	%ra, [%sp + 12]
"00111011110000010000000000000100",	-- 3032: 	lw	%r1, [%sp + 4]
"00111011110000100000000000001001",	-- 3033: 	lw	%r2, [%sp + 9]
"10000100010000010000100000000000",	-- 3034: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3035: 	lf	%f1, [%r1 + 0]
"00111111111111100000000000001100",	-- 3036: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3037: 	addi	%sp, %sp, 13
"01011000000000000000010011110011",	-- 3038: 	jal	fless.2532
"10101011110111100000000000001101",	-- 3039: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3040: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000000",	-- 3041: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3042: 	bneq	%r1, %r2, bneq_else.8990
"11001100000000010000000000000000",	-- 3043: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3044: 	jr	%ra
	-- bneq_else.8990:
"00111011110000010000000000000010",	-- 3045: 	lw	%r1, [%sp + 2]
"00111011110000100000000000000111",	-- 3046: 	lw	%r2, [%sp + 7]
"10000100010000010001000000000000",	-- 3047: 	add	%r2, %r2, %r1
"10010000010000000000000000000000",	-- 3048: 	lf	%f0, [%r2 + 0]
"10010011110000010000000000001011",	-- 3049: 	lf	%f1, [%sp + 11]
"11101000001000000000000000000000",	-- 3050: 	mulf	%f0, %f1, %f0
"10010011110000100000000000000001",	-- 3051: 	lf	%f2, [%sp + 1]
"11100000000000100000000000000000",	-- 3052: 	addf	%f0, %f0, %f2
"00111111111111100000000000001100",	-- 3053: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3054: 	addi	%sp, %sp, 13
"01011000000000000010101001001111",	-- 3055: 	jal	yj_fabs
"10101011110111100000000000001101",	-- 3056: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3057: 	lw	%ra, [%sp + 12]
"00111011110000010000000000000010",	-- 3058: 	lw	%r1, [%sp + 2]
"00111011110000100000000000001001",	-- 3059: 	lw	%r2, [%sp + 9]
"10000100010000010000100000000000",	-- 3060: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3061: 	lf	%f1, [%r1 + 0]
"00111111111111100000000000001100",	-- 3062: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3063: 	addi	%sp, %sp, 13
"01011000000000000000010011110011",	-- 3064: 	jal	fless.2532
"10101011110111100000000000001101",	-- 3065: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3066: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000000",	-- 3067: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3068: 	bneq	%r1, %r2, bneq_else.8991
"11001100000000010000000000000000",	-- 3069: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3070: 	jr	%ra
	-- bneq_else.8991:
"11001100000000010000000000000000",	-- 3071: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 3072: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3073: 	add	%r1, %r2, %r1
"10010011110000000000000000001011",	-- 3074: 	lf	%f0, [%sp + 11]
"10110000000000010000000000000000",	-- 3075: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 3076: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 3077: 	jr	%ra
	-- bneq_else.8989:
"11001100000000010000000000000000",	-- 3078: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3079: 	jr	%ra
	-- solver_rect.2725:
"00111011011110110000000000000001",	-- 3080: 	lw	%r27, [%r27 + 1]
"11001100000000110000000000000000",	-- 3081: 	lli	%r3, 0
"11001100000001000000000000000001",	-- 3082: 	lli	%r4, 1
"11001100000001010000000000000010",	-- 3083: 	lli	%r5, 2
"10110000000111100000000000000000",	-- 3084: 	sf	%f0, [%sp + 0]
"10110000010111100000000000000001",	-- 3085: 	sf	%f2, [%sp + 1]
"10110000001111100000000000000010",	-- 3086: 	sf	%f1, [%sp + 2]
"00111100010111100000000000000011",	-- 3087: 	sw	%r2, [%sp + 3]
"00111100001111100000000000000100",	-- 3088: 	sw	%r1, [%sp + 4]
"00111111011111100000000000000101",	-- 3089: 	sw	%r27, [%sp + 5]
"00111111111111100000000000000110",	-- 3090: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 3091: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 3092: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 3093: 	jalr	%r26
"10101011110111100000000000000111",	-- 3094: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 3095: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 3096: 	lli	%r2, 0
"00101000001000100000000000101001",	-- 3097: 	bneq	%r1, %r2, bneq_else.8992
"11001100000000110000000000000001",	-- 3098: 	lli	%r3, 1
"11001100000001000000000000000010",	-- 3099: 	lli	%r4, 2
"11001100000001010000000000000000",	-- 3100: 	lli	%r5, 0
"10010011110000000000000000000010",	-- 3101: 	lf	%f0, [%sp + 2]
"10010011110000010000000000000001",	-- 3102: 	lf	%f1, [%sp + 1]
"10010011110000100000000000000000",	-- 3103: 	lf	%f2, [%sp + 0]
"00111011110000010000000000000100",	-- 3104: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000011",	-- 3105: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000101",	-- 3106: 	lw	%r27, [%sp + 5]
"00111111111111100000000000000110",	-- 3107: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 3108: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 3109: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 3110: 	jalr	%r26
"10101011110111100000000000000111",	-- 3111: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 3112: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 3113: 	lli	%r2, 0
"00101000001000100000000000010110",	-- 3114: 	bneq	%r1, %r2, bneq_else.8993
"11001100000000110000000000000010",	-- 3115: 	lli	%r3, 2
"11001100000001000000000000000000",	-- 3116: 	lli	%r4, 0
"11001100000001010000000000000001",	-- 3117: 	lli	%r5, 1
"10010011110000000000000000000001",	-- 3118: 	lf	%f0, [%sp + 1]
"10010011110000010000000000000000",	-- 3119: 	lf	%f1, [%sp + 0]
"10010011110000100000000000000010",	-- 3120: 	lf	%f2, [%sp + 2]
"00111011110000010000000000000100",	-- 3121: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000011",	-- 3122: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000101",	-- 3123: 	lw	%r27, [%sp + 5]
"00111111111111100000000000000110",	-- 3124: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 3125: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 3126: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 3127: 	jalr	%r26
"10101011110111100000000000000111",	-- 3128: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 3129: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 3130: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3131: 	bneq	%r1, %r2, bneq_else.8994
"11001100000000010000000000000000",	-- 3132: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3133: 	jr	%ra
	-- bneq_else.8994:
"11001100000000010000000000000011",	-- 3134: 	lli	%r1, 3
"01001111111000000000000000000000",	-- 3135: 	jr	%ra
	-- bneq_else.8993:
"11001100000000010000000000000010",	-- 3136: 	lli	%r1, 2
"01001111111000000000000000000000",	-- 3137: 	jr	%ra
	-- bneq_else.8992:
"11001100000000010000000000000001",	-- 3138: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 3139: 	jr	%ra
	-- solver_surface.2731:
"00111011011000110000000000000001",	-- 3140: 	lw	%r3, [%r27 + 1]
"00111100011111100000000000000000",	-- 3141: 	sw	%r3, [%sp + 0]
"10110000010111100000000000000001",	-- 3142: 	sf	%f2, [%sp + 1]
"10110000001111100000000000000010",	-- 3143: 	sf	%f1, [%sp + 2]
"10110000000111100000000000000011",	-- 3144: 	sf	%f0, [%sp + 3]
"00111100010111100000000000000100",	-- 3145: 	sw	%r2, [%sp + 4]
"00111111111111100000000000000101",	-- 3146: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 3147: 	addi	%sp, %sp, 6
"01011000000000000000011001101001",	-- 3148: 	jal	o_param_abc.2638
"10101011110111100000000000000110",	-- 3149: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 3150: 	lw	%ra, [%sp + 5]
"10000100000000010001000000000000",	-- 3151: 	add	%r2, %r0, %r1
"00111011110000010000000000000100",	-- 3152: 	lw	%r1, [%sp + 4]
"00111100010111100000000000000101",	-- 3153: 	sw	%r2, [%sp + 5]
"00111111111111100000000000000110",	-- 3154: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 3155: 	addi	%sp, %sp, 7
"01011000000000000000010110100111",	-- 3156: 	jal	veciprod.2597
"10101011110111100000000000000111",	-- 3157: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 3158: 	lw	%ra, [%sp + 6]
"10110000000111100000000000000110",	-- 3159: 	sf	%f0, [%sp + 6]
"00111111111111100000000000000111",	-- 3160: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 3161: 	addi	%sp, %sp, 8
"01011000000000000000010011010110",	-- 3162: 	jal	fispos.2522
"10101011110111100000000000001000",	-- 3163: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 3164: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000000",	-- 3165: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3166: 	bneq	%r1, %r2, bneq_else.8995
"11001100000000010000000000000000",	-- 3167: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3168: 	jr	%ra
	-- bneq_else.8995:
"11001100000000010000000000000000",	-- 3169: 	lli	%r1, 0
"10010011110000000000000000000011",	-- 3170: 	lf	%f0, [%sp + 3]
"10010011110000010000000000000010",	-- 3171: 	lf	%f1, [%sp + 2]
"10010011110000100000000000000001",	-- 3172: 	lf	%f2, [%sp + 1]
"00111011110000100000000000000101",	-- 3173: 	lw	%r2, [%sp + 5]
"00111100001111100000000000000111",	-- 3174: 	sw	%r1, [%sp + 7]
"10000100000000100000100000000000",	-- 3175: 	add	%r1, %r0, %r2
"00111111111111100000000000001000",	-- 3176: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 3177: 	addi	%sp, %sp, 9
"01011000000000000000010110111111",	-- 3178: 	jal	veciprod2.2600
"10101011110111100000000000001001",	-- 3179: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 3180: 	lw	%ra, [%sp + 8]
"00111111111111100000000000001000",	-- 3181: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 3182: 	addi	%sp, %sp, 9
"01011000000000000010101001010001",	-- 3183: 	jal	yj_fneg
"10101011110111100000000000001001",	-- 3184: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 3185: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000110",	-- 3186: 	lf	%f1, [%sp + 6]
"11101100000000010000000000000000",	-- 3187: 	divf	%f0, %f0, %f1
"00111011110000010000000000000111",	-- 3188: 	lw	%r1, [%sp + 7]
"00111011110000100000000000000000",	-- 3189: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3190: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 3191: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 3192: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 3193: 	jr	%ra
	-- quadratic.2737:
"10110000000111100000000000000000",	-- 3194: 	sf	%f0, [%sp + 0]
"10110000010111100000000000000001",	-- 3195: 	sf	%f2, [%sp + 1]
"10110000001111100000000000000010",	-- 3196: 	sf	%f1, [%sp + 2]
"00111100001111100000000000000011",	-- 3197: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 3198: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 3199: 	addi	%sp, %sp, 5
"01011000000000000000010011110001",	-- 3200: 	jal	fsqr.2530
"10101011110111100000000000000101",	-- 3201: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 3202: 	lw	%ra, [%sp + 4]
"00111011110000010000000000000011",	-- 3203: 	lw	%r1, [%sp + 3]
"10110000000111100000000000000100",	-- 3204: 	sf	%f0, [%sp + 4]
"00111111111111100000000000000101",	-- 3205: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 3206: 	addi	%sp, %sp, 6
"01011000000000000000011001011010",	-- 3207: 	jal	o_param_a.2632
"10101011110111100000000000000110",	-- 3208: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 3209: 	lw	%ra, [%sp + 5]
"10010011110000010000000000000100",	-- 3210: 	lf	%f1, [%sp + 4]
"11101000001000000000000000000000",	-- 3211: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000010",	-- 3212: 	lf	%f1, [%sp + 2]
"10110000000111100000000000000101",	-- 3213: 	sf	%f0, [%sp + 5]
"00001100001000000000000000000000",	-- 3214: 	movf	%f0, %f1
"00111111111111100000000000000110",	-- 3215: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 3216: 	addi	%sp, %sp, 7
"01011000000000000000010011110001",	-- 3217: 	jal	fsqr.2530
"10101011110111100000000000000111",	-- 3218: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 3219: 	lw	%ra, [%sp + 6]
"00111011110000010000000000000011",	-- 3220: 	lw	%r1, [%sp + 3]
"10110000000111100000000000000110",	-- 3221: 	sf	%f0, [%sp + 6]
"00111111111111100000000000000111",	-- 3222: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 3223: 	addi	%sp, %sp, 8
"01011000000000000000011001011111",	-- 3224: 	jal	o_param_b.2634
"10101011110111100000000000001000",	-- 3225: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 3226: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000110",	-- 3227: 	lf	%f1, [%sp + 6]
"11101000001000000000000000000000",	-- 3228: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000101",	-- 3229: 	lf	%f1, [%sp + 5]
"11100000001000000000000000000000",	-- 3230: 	addf	%f0, %f1, %f0
"10010011110000010000000000000001",	-- 3231: 	lf	%f1, [%sp + 1]
"10110000000111100000000000000111",	-- 3232: 	sf	%f0, [%sp + 7]
"00001100001000000000000000000000",	-- 3233: 	movf	%f0, %f1
"00111111111111100000000000001000",	-- 3234: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 3235: 	addi	%sp, %sp, 9
"01011000000000000000010011110001",	-- 3236: 	jal	fsqr.2530
"10101011110111100000000000001001",	-- 3237: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 3238: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000011",	-- 3239: 	lw	%r1, [%sp + 3]
"10110000000111100000000000001000",	-- 3240: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 3241: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 3242: 	addi	%sp, %sp, 10
"01011000000000000000011001100100",	-- 3243: 	jal	o_param_c.2636
"10101011110111100000000000001010",	-- 3244: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 3245: 	lw	%ra, [%sp + 9]
"10010011110000010000000000001000",	-- 3246: 	lf	%f1, [%sp + 8]
"11101000001000000000000000000000",	-- 3247: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000111",	-- 3248: 	lf	%f1, [%sp + 7]
"11100000001000000000000000000000",	-- 3249: 	addf	%f0, %f1, %f0
"00111011110000010000000000000011",	-- 3250: 	lw	%r1, [%sp + 3]
"10110000000111100000000000001001",	-- 3251: 	sf	%f0, [%sp + 9]
"00111111111111100000000000001010",	-- 3252: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 3253: 	addi	%sp, %sp, 11
"01011000000000000000011001011000",	-- 3254: 	jal	o_isrot.2630
"10101011110111100000000000001011",	-- 3255: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 3256: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 3257: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3258: 	bneq	%r1, %r2, bneq_else.8996
"10010011110000000000000000001001",	-- 3259: 	lf	%f0, [%sp + 9]
"01001111111000000000000000000000",	-- 3260: 	jr	%ra
	-- bneq_else.8996:
"10010011110000000000000000000001",	-- 3261: 	lf	%f0, [%sp + 1]
"10010011110000010000000000000010",	-- 3262: 	lf	%f1, [%sp + 2]
"11101000001000000001000000000000",	-- 3263: 	mulf	%f2, %f1, %f0
"00111011110000010000000000000011",	-- 3264: 	lw	%r1, [%sp + 3]
"10110000010111100000000000001010",	-- 3265: 	sf	%f2, [%sp + 10]
"00111111111111100000000000001011",	-- 3266: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 3267: 	addi	%sp, %sp, 12
"01011000000000000000011010010011",	-- 3268: 	jal	o_param_r1.2656
"10101011110111100000000000001100",	-- 3269: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3270: 	lw	%ra, [%sp + 11]
"10010011110000010000000000001010",	-- 3271: 	lf	%f1, [%sp + 10]
"11101000001000000000000000000000",	-- 3272: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001001",	-- 3273: 	lf	%f1, [%sp + 9]
"11100000001000000000000000000000",	-- 3274: 	addf	%f0, %f1, %f0
"10010011110000010000000000000000",	-- 3275: 	lf	%f1, [%sp + 0]
"10010011110000100000000000000001",	-- 3276: 	lf	%f2, [%sp + 1]
"11101000010000010001000000000000",	-- 3277: 	mulf	%f2, %f2, %f1
"00111011110000010000000000000011",	-- 3278: 	lw	%r1, [%sp + 3]
"10110000000111100000000000001011",	-- 3279: 	sf	%f0, [%sp + 11]
"10110000010111100000000000001100",	-- 3280: 	sf	%f2, [%sp + 12]
"00111111111111100000000000001101",	-- 3281: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 3282: 	addi	%sp, %sp, 14
"01011000000000000000011010011000",	-- 3283: 	jal	o_param_r2.2658
"10101011110111100000000000001110",	-- 3284: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 3285: 	lw	%ra, [%sp + 13]
"10010011110000010000000000001100",	-- 3286: 	lf	%f1, [%sp + 12]
"11101000001000000000000000000000",	-- 3287: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001011",	-- 3288: 	lf	%f1, [%sp + 11]
"11100000001000000000000000000000",	-- 3289: 	addf	%f0, %f1, %f0
"10010011110000010000000000000010",	-- 3290: 	lf	%f1, [%sp + 2]
"10010011110000100000000000000000",	-- 3291: 	lf	%f2, [%sp + 0]
"11101000010000010000100000000000",	-- 3292: 	mulf	%f1, %f2, %f1
"00111011110000010000000000000011",	-- 3293: 	lw	%r1, [%sp + 3]
"10110000000111100000000000001101",	-- 3294: 	sf	%f0, [%sp + 13]
"10110000001111100000000000001110",	-- 3295: 	sf	%f1, [%sp + 14]
"00111111111111100000000000001111",	-- 3296: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 3297: 	addi	%sp, %sp, 16
"01011000000000000000011010011101",	-- 3298: 	jal	o_param_r3.2660
"10101011110111100000000000010000",	-- 3299: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 3300: 	lw	%ra, [%sp + 15]
"10010011110000010000000000001110",	-- 3301: 	lf	%f1, [%sp + 14]
"11101000001000000000000000000000",	-- 3302: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001101",	-- 3303: 	lf	%f1, [%sp + 13]
"11100000001000000000000000000000",	-- 3304: 	addf	%f0, %f1, %f0
"01001111111000000000000000000000",	-- 3305: 	jr	%ra
	-- bilinear.2742:
"11101000000000110011000000000000",	-- 3306: 	mulf	%f6, %f0, %f3
"10110000011111100000000000000000",	-- 3307: 	sf	%f3, [%sp + 0]
"10110000000111100000000000000001",	-- 3308: 	sf	%f0, [%sp + 1]
"10110000101111100000000000000010",	-- 3309: 	sf	%f5, [%sp + 2]
"10110000010111100000000000000011",	-- 3310: 	sf	%f2, [%sp + 3]
"00111100001111100000000000000100",	-- 3311: 	sw	%r1, [%sp + 4]
"10110000100111100000000000000101",	-- 3312: 	sf	%f4, [%sp + 5]
"10110000001111100000000000000110",	-- 3313: 	sf	%f1, [%sp + 6]
"10110000110111100000000000000111",	-- 3314: 	sf	%f6, [%sp + 7]
"00111111111111100000000000001000",	-- 3315: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 3316: 	addi	%sp, %sp, 9
"01011000000000000000011001011010",	-- 3317: 	jal	o_param_a.2632
"10101011110111100000000000001001",	-- 3318: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 3319: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000111",	-- 3320: 	lf	%f1, [%sp + 7]
"11101000001000000000000000000000",	-- 3321: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000101",	-- 3322: 	lf	%f1, [%sp + 5]
"10010011110000100000000000000110",	-- 3323: 	lf	%f2, [%sp + 6]
"11101000010000010001100000000000",	-- 3324: 	mulf	%f3, %f2, %f1
"00111011110000010000000000000100",	-- 3325: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001000",	-- 3326: 	sf	%f0, [%sp + 8]
"10110000011111100000000000001001",	-- 3327: 	sf	%f3, [%sp + 9]
"00111111111111100000000000001010",	-- 3328: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 3329: 	addi	%sp, %sp, 11
"01011000000000000000011001011111",	-- 3330: 	jal	o_param_b.2634
"10101011110111100000000000001011",	-- 3331: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 3332: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 3333: 	lf	%f1, [%sp + 9]
"11101000001000000000000000000000",	-- 3334: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001000",	-- 3335: 	lf	%f1, [%sp + 8]
"11100000001000000000000000000000",	-- 3336: 	addf	%f0, %f1, %f0
"10010011110000010000000000000010",	-- 3337: 	lf	%f1, [%sp + 2]
"10010011110000100000000000000011",	-- 3338: 	lf	%f2, [%sp + 3]
"11101000010000010001100000000000",	-- 3339: 	mulf	%f3, %f2, %f1
"00111011110000010000000000000100",	-- 3340: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001010",	-- 3341: 	sf	%f0, [%sp + 10]
"10110000011111100000000000001011",	-- 3342: 	sf	%f3, [%sp + 11]
"00111111111111100000000000001100",	-- 3343: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3344: 	addi	%sp, %sp, 13
"01011000000000000000011001100100",	-- 3345: 	jal	o_param_c.2636
"10101011110111100000000000001101",	-- 3346: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3347: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001011",	-- 3348: 	lf	%f1, [%sp + 11]
"11101000001000000000000000000000",	-- 3349: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001010",	-- 3350: 	lf	%f1, [%sp + 10]
"11100000001000000000000000000000",	-- 3351: 	addf	%f0, %f1, %f0
"00111011110000010000000000000100",	-- 3352: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001100",	-- 3353: 	sf	%f0, [%sp + 12]
"00111111111111100000000000001101",	-- 3354: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 3355: 	addi	%sp, %sp, 14
"01011000000000000000011001011000",	-- 3356: 	jal	o_isrot.2630
"10101011110111100000000000001110",	-- 3357: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 3358: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 3359: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3360: 	bneq	%r1, %r2, bneq_else.8997
"10010011110000000000000000001100",	-- 3361: 	lf	%f0, [%sp + 12]
"01001111111000000000000000000000",	-- 3362: 	jr	%ra
	-- bneq_else.8997:
"10010011110000000000000000000101",	-- 3363: 	lf	%f0, [%sp + 5]
"10010011110000010000000000000011",	-- 3364: 	lf	%f1, [%sp + 3]
"11101000001000000001000000000000",	-- 3365: 	mulf	%f2, %f1, %f0
"10010011110000110000000000000010",	-- 3366: 	lf	%f3, [%sp + 2]
"10010011110001000000000000000110",	-- 3367: 	lf	%f4, [%sp + 6]
"11101000100000110010100000000000",	-- 3368: 	mulf	%f5, %f4, %f3
"11100000010001010001000000000000",	-- 3369: 	addf	%f2, %f2, %f5
"00111011110000010000000000000100",	-- 3370: 	lw	%r1, [%sp + 4]
"10110000010111100000000000001101",	-- 3371: 	sf	%f2, [%sp + 13]
"00111111111111100000000000001110",	-- 3372: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 3373: 	addi	%sp, %sp, 15
"01011000000000000000011010010011",	-- 3374: 	jal	o_param_r1.2656
"10101011110111100000000000001111",	-- 3375: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 3376: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001101",	-- 3377: 	lf	%f1, [%sp + 13]
"11101000001000000000000000000000",	-- 3378: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000010",	-- 3379: 	lf	%f1, [%sp + 2]
"10010011110000100000000000000001",	-- 3380: 	lf	%f2, [%sp + 1]
"11101000010000010000100000000000",	-- 3381: 	mulf	%f1, %f2, %f1
"10010011110000110000000000000000",	-- 3382: 	lf	%f3, [%sp + 0]
"10010011110001000000000000000011",	-- 3383: 	lf	%f4, [%sp + 3]
"11101000100000110010000000000000",	-- 3384: 	mulf	%f4, %f4, %f3
"11100000001001000000100000000000",	-- 3385: 	addf	%f1, %f1, %f4
"00111011110000010000000000000100",	-- 3386: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001110",	-- 3387: 	sf	%f0, [%sp + 14]
"10110000001111100000000000001111",	-- 3388: 	sf	%f1, [%sp + 15]
"00111111111111100000000000010000",	-- 3389: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 3390: 	addi	%sp, %sp, 17
"01011000000000000000011010011000",	-- 3391: 	jal	o_param_r2.2658
"10101011110111100000000000010001",	-- 3392: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 3393: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001111",	-- 3394: 	lf	%f1, [%sp + 15]
"11101000001000000000000000000000",	-- 3395: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001110",	-- 3396: 	lf	%f1, [%sp + 14]
"11100000001000000000000000000000",	-- 3397: 	addf	%f0, %f1, %f0
"10010011110000010000000000000101",	-- 3398: 	lf	%f1, [%sp + 5]
"10010011110000100000000000000001",	-- 3399: 	lf	%f2, [%sp + 1]
"11101000010000010000100000000000",	-- 3400: 	mulf	%f1, %f2, %f1
"10010011110000100000000000000000",	-- 3401: 	lf	%f2, [%sp + 0]
"10010011110000110000000000000110",	-- 3402: 	lf	%f3, [%sp + 6]
"11101000011000100001000000000000",	-- 3403: 	mulf	%f2, %f3, %f2
"11100000001000100000100000000000",	-- 3404: 	addf	%f1, %f1, %f2
"00111011110000010000000000000100",	-- 3405: 	lw	%r1, [%sp + 4]
"10110000000111100000000000010000",	-- 3406: 	sf	%f0, [%sp + 16]
"10110000001111100000000000010001",	-- 3407: 	sf	%f1, [%sp + 17]
"00111111111111100000000000010010",	-- 3408: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 3409: 	addi	%sp, %sp, 19
"01011000000000000000011010011101",	-- 3410: 	jal	o_param_r3.2660
"10101011110111100000000000010011",	-- 3411: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 3412: 	lw	%ra, [%sp + 18]
"10010011110000010000000000010001",	-- 3413: 	lf	%f1, [%sp + 17]
"11101000001000000000000000000000",	-- 3414: 	mulf	%f0, %f1, %f0
"10010011110000010000000000010000",	-- 3415: 	lf	%f1, [%sp + 16]
"11100000001000000000000000000000",	-- 3416: 	addf	%f0, %f1, %f0
"00111111111111100000000000010010",	-- 3417: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 3418: 	addi	%sp, %sp, 19
"01011000000000000000010011101101",	-- 3419: 	jal	fhalf.2528
"10101011110111100000000000010011",	-- 3420: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 3421: 	lw	%ra, [%sp + 18]
"10010011110000010000000000001100",	-- 3422: 	lf	%f1, [%sp + 12]
"11100000001000000000000000000000",	-- 3423: 	addf	%f0, %f1, %f0
"01001111111000000000000000000000",	-- 3424: 	jr	%ra
	-- solver_second.2750:
"00111011011000110000000000000001",	-- 3425: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 3426: 	lli	%r4, 0
"10000100010001000010000000000000",	-- 3427: 	add	%r4, %r2, %r4
"10010000100000110000000000000000",	-- 3428: 	lf	%f3, [%r4 + 0]
"11001100000001000000000000000001",	-- 3429: 	lli	%r4, 1
"10000100010001000010000000000000",	-- 3430: 	add	%r4, %r2, %r4
"10010000100001000000000000000000",	-- 3431: 	lf	%f4, [%r4 + 0]
"11001100000001000000000000000010",	-- 3432: 	lli	%r4, 2
"10000100010001000010000000000000",	-- 3433: 	add	%r4, %r2, %r4
"10010000100001010000000000000000",	-- 3434: 	lf	%f5, [%r4 + 0]
"00111100011111100000000000000000",	-- 3435: 	sw	%r3, [%sp + 0]
"10110000010111100000000000000001",	-- 3436: 	sf	%f2, [%sp + 1]
"10110000001111100000000000000010",	-- 3437: 	sf	%f1, [%sp + 2]
"10110000000111100000000000000011",	-- 3438: 	sf	%f0, [%sp + 3]
"00111100001111100000000000000100",	-- 3439: 	sw	%r1, [%sp + 4]
"00111100010111100000000000000101",	-- 3440: 	sw	%r2, [%sp + 5]
"00001100101000100000000000000000",	-- 3441: 	movf	%f2, %f5
"00001100100000010000000000000000",	-- 3442: 	movf	%f1, %f4
"00001100011000000000000000000000",	-- 3443: 	movf	%f0, %f3
"00111111111111100000000000000110",	-- 3444: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 3445: 	addi	%sp, %sp, 7
"01011000000000000000110001111010",	-- 3446: 	jal	quadratic.2737
"10101011110111100000000000000111",	-- 3447: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 3448: 	lw	%ra, [%sp + 6]
"10110000000111100000000000000110",	-- 3449: 	sf	%f0, [%sp + 6]
"00111111111111100000000000000111",	-- 3450: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 3451: 	addi	%sp, %sp, 8
"01011000000000000000010011100100",	-- 3452: 	jal	fiszero.2526
"10101011110111100000000000001000",	-- 3453: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 3454: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000000",	-- 3455: 	lli	%r2, 0
"00101000001000100000000001100111",	-- 3456: 	bneq	%r1, %r2, bneq_else.8998
"11001100000000010000000000000000",	-- 3457: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 3458: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 3459: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3460: 	lf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 3461: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 3462: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3463: 	lf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 3464: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 3465: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 3466: 	lf	%f2, [%r1 + 0]
"10010011110000110000000000000011",	-- 3467: 	lf	%f3, [%sp + 3]
"10010011110001000000000000000010",	-- 3468: 	lf	%f4, [%sp + 2]
"10010011110001010000000000000001",	-- 3469: 	lf	%f5, [%sp + 1]
"00111011110000010000000000000100",	-- 3470: 	lw	%r1, [%sp + 4]
"00111111111111100000000000000111",	-- 3471: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 3472: 	addi	%sp, %sp, 8
"01011000000000000000110011101010",	-- 3473: 	jal	bilinear.2742
"10101011110111100000000000001000",	-- 3474: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 3475: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000011",	-- 3476: 	lf	%f1, [%sp + 3]
"10010011110000100000000000000010",	-- 3477: 	lf	%f2, [%sp + 2]
"10010011110000110000000000000001",	-- 3478: 	lf	%f3, [%sp + 1]
"00111011110000010000000000000100",	-- 3479: 	lw	%r1, [%sp + 4]
"10110000000111100000000000000111",	-- 3480: 	sf	%f0, [%sp + 7]
"00001100001000000000000000000000",	-- 3481: 	movf	%f0, %f1
"00001100010000010000000000000000",	-- 3482: 	movf	%f1, %f2
"00001100011000100000000000000000",	-- 3483: 	movf	%f2, %f3
"00111111111111100000000000001000",	-- 3484: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 3485: 	addi	%sp, %sp, 9
"01011000000000000000110001111010",	-- 3486: 	jal	quadratic.2737
"10101011110111100000000000001001",	-- 3487: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 3488: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000100",	-- 3489: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001000",	-- 3490: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 3491: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 3492: 	addi	%sp, %sp, 10
"01011000000000000000011001010010",	-- 3493: 	jal	o_form.2624
"10101011110111100000000000001010",	-- 3494: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 3495: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000011",	-- 3496: 	lli	%r2, 3
"00101000001000100000000000000110",	-- 3497: 	bneq	%r1, %r2, bneq_else.8999
"00010100000000000000000000000000",	-- 3498: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 3499: 	lhif	%f0, 1.000000
"10010011110000010000000000001000",	-- 3500: 	lf	%f1, [%sp + 8]
"11100100001000000000000000000000",	-- 3501: 	subf	%f0, %f1, %f0
"01010100000000000000110110110000",	-- 3502: 	j	bneq_cont.9000
	-- bneq_else.8999:
"10010011110000000000000000001000",	-- 3503: 	lf	%f0, [%sp + 8]
	-- bneq_cont.9000:
"10010011110000010000000000000111",	-- 3504: 	lf	%f1, [%sp + 7]
"10110000000111100000000000001001",	-- 3505: 	sf	%f0, [%sp + 9]
"00001100001000000000000000000000",	-- 3506: 	movf	%f0, %f1
"00111111111111100000000000001010",	-- 3507: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 3508: 	addi	%sp, %sp, 11
"01011000000000000000010011110001",	-- 3509: 	jal	fsqr.2530
"10101011110111100000000000001011",	-- 3510: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 3511: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 3512: 	lf	%f1, [%sp + 9]
"10010011110000100000000000000110",	-- 3513: 	lf	%f2, [%sp + 6]
"11101000010000010000100000000000",	-- 3514: 	mulf	%f1, %f2, %f1
"11100100000000010000000000000000",	-- 3515: 	subf	%f0, %f0, %f1
"10110000000111100000000000001010",	-- 3516: 	sf	%f0, [%sp + 10]
"00111111111111100000000000001011",	-- 3517: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 3518: 	addi	%sp, %sp, 12
"01011000000000000000010011010110",	-- 3519: 	jal	fispos.2522
"10101011110111100000000000001100",	-- 3520: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3521: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 3522: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3523: 	bneq	%r1, %r2, bneq_else.9001
"11001100000000010000000000000000",	-- 3524: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3525: 	jr	%ra
	-- bneq_else.9001:
"10010011110000000000000000001010",	-- 3526: 	lf	%f0, [%sp + 10]
"00111111111111100000000000001011",	-- 3527: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 3528: 	addi	%sp, %sp, 12
"01011000000000000010101000110000",	-- 3529: 	jal	yj_sqrt
"10101011110111100000000000001100",	-- 3530: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3531: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000100",	-- 3532: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001011",	-- 3533: 	sf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 3534: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3535: 	addi	%sp, %sp, 13
"01011000000000000000011001010110",	-- 3536: 	jal	o_isinvert.2628
"10101011110111100000000000001101",	-- 3537: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3538: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000000",	-- 3539: 	lli	%r2, 0
"00101000001000100000000000001000",	-- 3540: 	bneq	%r1, %r2, bneq_else.9002
"10010011110000000000000000001011",	-- 3541: 	lf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 3542: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3543: 	addi	%sp, %sp, 13
"01011000000000000010101001010001",	-- 3544: 	jal	yj_fneg
"10101011110111100000000000001101",	-- 3545: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3546: 	lw	%ra, [%sp + 12]
"01010100000000000000110111011101",	-- 3547: 	j	bneq_cont.9003
	-- bneq_else.9002:
"10010011110000000000000000001011",	-- 3548: 	lf	%f0, [%sp + 11]
	-- bneq_cont.9003:
"11001100000000010000000000000000",	-- 3549: 	lli	%r1, 0
"10010011110000010000000000000111",	-- 3550: 	lf	%f1, [%sp + 7]
"11100100000000010000000000000000",	-- 3551: 	subf	%f0, %f0, %f1
"10010011110000010000000000000110",	-- 3552: 	lf	%f1, [%sp + 6]
"11101100000000010000000000000000",	-- 3553: 	divf	%f0, %f0, %f1
"00111011110000100000000000000000",	-- 3554: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3555: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 3556: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 3557: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 3558: 	jr	%ra
	-- bneq_else.8998:
"11001100000000010000000000000000",	-- 3559: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3560: 	jr	%ra
	-- solver.2756:
"00111011011001000000000000000100",	-- 3561: 	lw	%r4, [%r27 + 4]
"00111011011001010000000000000011",	-- 3562: 	lw	%r5, [%r27 + 3]
"00111011011001100000000000000010",	-- 3563: 	lw	%r6, [%r27 + 2]
"00111011011001110000000000000001",	-- 3564: 	lw	%r7, [%r27 + 1]
"10000100111000010000100000000000",	-- 3565: 	add	%r1, %r7, %r1
"00111000001000010000000000000000",	-- 3566: 	lw	%r1, [%r1 + 0]
"11001100000001110000000000000000",	-- 3567: 	lli	%r7, 0
"10000100011001110011100000000000",	-- 3568: 	add	%r7, %r3, %r7
"10010000111000000000000000000000",	-- 3569: 	lf	%f0, [%r7 + 0]
"00111100101111100000000000000000",	-- 3570: 	sw	%r5, [%sp + 0]
"00111100100111100000000000000001",	-- 3571: 	sw	%r4, [%sp + 1]
"00111100010111100000000000000010",	-- 3572: 	sw	%r2, [%sp + 2]
"00111100110111100000000000000011",	-- 3573: 	sw	%r6, [%sp + 3]
"00111100001111100000000000000100",	-- 3574: 	sw	%r1, [%sp + 4]
"00111100011111100000000000000101",	-- 3575: 	sw	%r3, [%sp + 5]
"10110000000111100000000000000110",	-- 3576: 	sf	%f0, [%sp + 6]
"00111111111111100000000000000111",	-- 3577: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 3578: 	addi	%sp, %sp, 8
"01011000000000000000011001101011",	-- 3579: 	jal	o_param_x.2640
"10101011110111100000000000001000",	-- 3580: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 3581: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000110",	-- 3582: 	lf	%f1, [%sp + 6]
"11100100001000000000000000000000",	-- 3583: 	subf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 3584: 	lli	%r1, 1
"00111011110000100000000000000101",	-- 3585: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 3586: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3587: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000100",	-- 3588: 	lw	%r1, [%sp + 4]
"10110000000111100000000000000111",	-- 3589: 	sf	%f0, [%sp + 7]
"10110000001111100000000000001000",	-- 3590: 	sf	%f1, [%sp + 8]
"00111111111111100000000000001001",	-- 3591: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 3592: 	addi	%sp, %sp, 10
"01011000000000000000011001110000",	-- 3593: 	jal	o_param_y.2642
"10101011110111100000000000001010",	-- 3594: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 3595: 	lw	%ra, [%sp + 9]
"10010011110000010000000000001000",	-- 3596: 	lf	%f1, [%sp + 8]
"11100100001000000000000000000000",	-- 3597: 	subf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 3598: 	lli	%r1, 2
"00111011110000100000000000000101",	-- 3599: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 3600: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3601: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000100",	-- 3602: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001001",	-- 3603: 	sf	%f0, [%sp + 9]
"10110000001111100000000000001010",	-- 3604: 	sf	%f1, [%sp + 10]
"00111111111111100000000000001011",	-- 3605: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 3606: 	addi	%sp, %sp, 12
"01011000000000000000011001110101",	-- 3607: 	jal	o_param_z.2644
"10101011110111100000000000001100",	-- 3608: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3609: 	lw	%ra, [%sp + 11]
"10010011110000010000000000001010",	-- 3610: 	lf	%f1, [%sp + 10]
"11100100001000000000000000000000",	-- 3611: 	subf	%f0, %f1, %f0
"00111011110000010000000000000100",	-- 3612: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001011",	-- 3613: 	sf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 3614: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3615: 	addi	%sp, %sp, 13
"01011000000000000000011001010010",	-- 3616: 	jal	o_form.2624
"10101011110111100000000000001101",	-- 3617: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3618: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000001",	-- 3619: 	lli	%r2, 1
"00101000001000100000000000001001",	-- 3620: 	bneq	%r1, %r2, bneq_else.9004
"10010011110000000000000000000111",	-- 3621: 	lf	%f0, [%sp + 7]
"10010011110000010000000000001001",	-- 3622: 	lf	%f1, [%sp + 9]
"10010011110000100000000000001011",	-- 3623: 	lf	%f2, [%sp + 11]
"00111011110000010000000000000100",	-- 3624: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000010",	-- 3625: 	lw	%r2, [%sp + 2]
"00111011110110110000000000000011",	-- 3626: 	lw	%r27, [%sp + 3]
"00111011011110100000000000000000",	-- 3627: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 3628: 	jr	%r26
	-- bneq_else.9004:
"11001100000000100000000000000010",	-- 3629: 	lli	%r2, 2
"00101000001000100000000000001001",	-- 3630: 	bneq	%r1, %r2, bneq_else.9005
"10010011110000000000000000000111",	-- 3631: 	lf	%f0, [%sp + 7]
"10010011110000010000000000001001",	-- 3632: 	lf	%f1, [%sp + 9]
"10010011110000100000000000001011",	-- 3633: 	lf	%f2, [%sp + 11]
"00111011110000010000000000000100",	-- 3634: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000010",	-- 3635: 	lw	%r2, [%sp + 2]
"00111011110110110000000000000001",	-- 3636: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 3637: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 3638: 	jr	%r26
	-- bneq_else.9005:
"10010011110000000000000000000111",	-- 3639: 	lf	%f0, [%sp + 7]
"10010011110000010000000000001001",	-- 3640: 	lf	%f1, [%sp + 9]
"10010011110000100000000000001011",	-- 3641: 	lf	%f2, [%sp + 11]
"00111011110000010000000000000100",	-- 3642: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000010",	-- 3643: 	lw	%r2, [%sp + 2]
"00111011110110110000000000000000",	-- 3644: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 3645: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 3646: 	jr	%r26
	-- solver_rect_fast.2760:
"00111011011001000000000000000001",	-- 3647: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 3648: 	lli	%r5, 0
"10000100011001010010100000000000",	-- 3649: 	add	%r5, %r3, %r5
"10010000101000110000000000000000",	-- 3650: 	lf	%f3, [%r5 + 0]
"11100100011000000001100000000000",	-- 3651: 	subf	%f3, %f3, %f0
"11001100000001010000000000000001",	-- 3652: 	lli	%r5, 1
"10000100011001010010100000000000",	-- 3653: 	add	%r5, %r3, %r5
"10010000101001000000000000000000",	-- 3654: 	lf	%f4, [%r5 + 0]
"11101000011001000001100000000000",	-- 3655: 	mulf	%f3, %f3, %f4
"11001100000001010000000000000001",	-- 3656: 	lli	%r5, 1
"10000100010001010010100000000000",	-- 3657: 	add	%r5, %r2, %r5
"10010000101001000000000000000000",	-- 3658: 	lf	%f4, [%r5 + 0]
"11101000011001000010000000000000",	-- 3659: 	mulf	%f4, %f3, %f4
"11100000100000010010000000000000",	-- 3660: 	addf	%f4, %f4, %f1
"00111100100111100000000000000000",	-- 3661: 	sw	%r4, [%sp + 0]
"10110000000111100000000000000001",	-- 3662: 	sf	%f0, [%sp + 1]
"10110000001111100000000000000010",	-- 3663: 	sf	%f1, [%sp + 2]
"00111100011111100000000000000011",	-- 3664: 	sw	%r3, [%sp + 3]
"10110000010111100000000000000100",	-- 3665: 	sf	%f2, [%sp + 4]
"10110000011111100000000000000101",	-- 3666: 	sf	%f3, [%sp + 5]
"00111100010111100000000000000110",	-- 3667: 	sw	%r2, [%sp + 6]
"00111100001111100000000000000111",	-- 3668: 	sw	%r1, [%sp + 7]
"00001100100000000000000000000000",	-- 3669: 	movf	%f0, %f4
"00111111111111100000000000001000",	-- 3670: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 3671: 	addi	%sp, %sp, 9
"01011000000000000010101001001111",	-- 3672: 	jal	yj_fabs
"10101011110111100000000000001001",	-- 3673: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 3674: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000111",	-- 3675: 	lw	%r1, [%sp + 7]
"10110000000111100000000000001000",	-- 3676: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 3677: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 3678: 	addi	%sp, %sp, 10
"01011000000000000000011001011111",	-- 3679: 	jal	o_param_b.2634
"10101011110111100000000000001010",	-- 3680: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 3681: 	lw	%ra, [%sp + 9]
"00001100000000010000000000000000",	-- 3682: 	movf	%f1, %f0
"10010011110000000000000000001000",	-- 3683: 	lf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 3684: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 3685: 	addi	%sp, %sp, 10
"01011000000000000000010011110011",	-- 3686: 	jal	fless.2532
"10101011110111100000000000001010",	-- 3687: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 3688: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000000",	-- 3689: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3690: 	bneq	%r1, %r2, bneq_else.9006
"11001100000000010000000000000000",	-- 3691: 	lli	%r1, 0
"01010100000000000000111010011010",	-- 3692: 	j	bneq_cont.9007
	-- bneq_else.9006:
"11001100000000010000000000000010",	-- 3693: 	lli	%r1, 2
"00111011110000100000000000000110",	-- 3694: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 3695: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3696: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000000101",	-- 3697: 	lf	%f1, [%sp + 5]
"11101000001000000000000000000000",	-- 3698: 	mulf	%f0, %f1, %f0
"10010011110000100000000000000100",	-- 3699: 	lf	%f2, [%sp + 4]
"11100000000000100000000000000000",	-- 3700: 	addf	%f0, %f0, %f2
"00111111111111100000000000001001",	-- 3701: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 3702: 	addi	%sp, %sp, 10
"01011000000000000010101001001111",	-- 3703: 	jal	yj_fabs
"10101011110111100000000000001010",	-- 3704: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 3705: 	lw	%ra, [%sp + 9]
"00111011110000010000000000000111",	-- 3706: 	lw	%r1, [%sp + 7]
"10110000000111100000000000001001",	-- 3707: 	sf	%f0, [%sp + 9]
"00111111111111100000000000001010",	-- 3708: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 3709: 	addi	%sp, %sp, 11
"01011000000000000000011001100100",	-- 3710: 	jal	o_param_c.2636
"10101011110111100000000000001011",	-- 3711: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 3712: 	lw	%ra, [%sp + 10]
"00001100000000010000000000000000",	-- 3713: 	movf	%f1, %f0
"10010011110000000000000000001001",	-- 3714: 	lf	%f0, [%sp + 9]
"00111111111111100000000000001010",	-- 3715: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 3716: 	addi	%sp, %sp, 11
"01011000000000000000010011110011",	-- 3717: 	jal	fless.2532
"10101011110111100000000000001011",	-- 3718: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 3719: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 3720: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3721: 	bneq	%r1, %r2, bneq_else.9008
"11001100000000010000000000000000",	-- 3722: 	lli	%r1, 0
"01010100000000000000111010011010",	-- 3723: 	j	bneq_cont.9009
	-- bneq_else.9008:
"11001100000000010000000000000001",	-- 3724: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 3725: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 3726: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3727: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000001010",	-- 3728: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 3729: 	addi	%sp, %sp, 11
"01011000000000000000010011100100",	-- 3730: 	jal	fiszero.2526
"10101011110111100000000000001011",	-- 3731: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 3732: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 3733: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3734: 	bneq	%r1, %r2, bneq_else.9010
"11001100000000010000000000000001",	-- 3735: 	lli	%r1, 1
"01010100000000000000111010011010",	-- 3736: 	j	bneq_cont.9011
	-- bneq_else.9010:
"11001100000000010000000000000000",	-- 3737: 	lli	%r1, 0
	-- bneq_cont.9011:
	-- bneq_cont.9009:
	-- bneq_cont.9007:
"11001100000000100000000000000000",	-- 3738: 	lli	%r2, 0
"00101000001000100000000011000011",	-- 3739: 	bneq	%r1, %r2, bneq_else.9012
"11001100000000010000000000000010",	-- 3740: 	lli	%r1, 2
"00111011110000100000000000000011",	-- 3741: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 3742: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3743: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000000010",	-- 3744: 	lf	%f1, [%sp + 2]
"11100100000000010000000000000000",	-- 3745: 	subf	%f0, %f0, %f1
"11001100000000010000000000000011",	-- 3746: 	lli	%r1, 3
"10000100010000010000100000000000",	-- 3747: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 3748: 	lf	%f2, [%r1 + 0]
"11101000000000100000000000000000",	-- 3749: 	mulf	%f0, %f0, %f2
"11001100000000010000000000000000",	-- 3750: 	lli	%r1, 0
"00111011110000110000000000000110",	-- 3751: 	lw	%r3, [%sp + 6]
"10000100011000010000100000000000",	-- 3752: 	add	%r1, %r3, %r1
"10010000001000100000000000000000",	-- 3753: 	lf	%f2, [%r1 + 0]
"11101000000000100001000000000000",	-- 3754: 	mulf	%f2, %f0, %f2
"10010011110000110000000000000001",	-- 3755: 	lf	%f3, [%sp + 1]
"11100000010000110001000000000000",	-- 3756: 	addf	%f2, %f2, %f3
"10110000000111100000000000001010",	-- 3757: 	sf	%f0, [%sp + 10]
"00001100010000000000000000000000",	-- 3758: 	movf	%f0, %f2
"00111111111111100000000000001011",	-- 3759: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 3760: 	addi	%sp, %sp, 12
"01011000000000000010101001001111",	-- 3761: 	jal	yj_fabs
"10101011110111100000000000001100",	-- 3762: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 3763: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000111",	-- 3764: 	lw	%r1, [%sp + 7]
"10110000000111100000000000001011",	-- 3765: 	sf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 3766: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3767: 	addi	%sp, %sp, 13
"01011000000000000000011001011010",	-- 3768: 	jal	o_param_a.2632
"10101011110111100000000000001101",	-- 3769: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3770: 	lw	%ra, [%sp + 12]
"00001100000000010000000000000000",	-- 3771: 	movf	%f1, %f0
"10010011110000000000000000001011",	-- 3772: 	lf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 3773: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3774: 	addi	%sp, %sp, 13
"01011000000000000000010011110011",	-- 3775: 	jal	fless.2532
"10101011110111100000000000001101",	-- 3776: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3777: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000000",	-- 3778: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3779: 	bneq	%r1, %r2, bneq_else.9013
"11001100000000010000000000000000",	-- 3780: 	lli	%r1, 0
"01010100000000000000111011110011",	-- 3781: 	j	bneq_cont.9014
	-- bneq_else.9013:
"11001100000000010000000000000010",	-- 3782: 	lli	%r1, 2
"00111011110000100000000000000110",	-- 3783: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 3784: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3785: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000001010",	-- 3786: 	lf	%f1, [%sp + 10]
"11101000001000000000000000000000",	-- 3787: 	mulf	%f0, %f1, %f0
"10010011110000100000000000000100",	-- 3788: 	lf	%f2, [%sp + 4]
"11100000000000100000000000000000",	-- 3789: 	addf	%f0, %f0, %f2
"00111111111111100000000000001100",	-- 3790: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 3791: 	addi	%sp, %sp, 13
"01011000000000000010101001001111",	-- 3792: 	jal	yj_fabs
"10101011110111100000000000001101",	-- 3793: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 3794: 	lw	%ra, [%sp + 12]
"00111011110000010000000000000111",	-- 3795: 	lw	%r1, [%sp + 7]
"10110000000111100000000000001100",	-- 3796: 	sf	%f0, [%sp + 12]
"00111111111111100000000000001101",	-- 3797: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 3798: 	addi	%sp, %sp, 14
"01011000000000000000011001100100",	-- 3799: 	jal	o_param_c.2636
"10101011110111100000000000001110",	-- 3800: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 3801: 	lw	%ra, [%sp + 13]
"00001100000000010000000000000000",	-- 3802: 	movf	%f1, %f0
"10010011110000000000000000001100",	-- 3803: 	lf	%f0, [%sp + 12]
"00111111111111100000000000001101",	-- 3804: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 3805: 	addi	%sp, %sp, 14
"01011000000000000000010011110011",	-- 3806: 	jal	fless.2532
"10101011110111100000000000001110",	-- 3807: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 3808: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 3809: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3810: 	bneq	%r1, %r2, bneq_else.9015
"11001100000000010000000000000000",	-- 3811: 	lli	%r1, 0
"01010100000000000000111011110011",	-- 3812: 	j	bneq_cont.9016
	-- bneq_else.9015:
"11001100000000010000000000000011",	-- 3813: 	lli	%r1, 3
"00111011110000100000000000000011",	-- 3814: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 3815: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3816: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000001101",	-- 3817: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 3818: 	addi	%sp, %sp, 14
"01011000000000000000010011100100",	-- 3819: 	jal	fiszero.2526
"10101011110111100000000000001110",	-- 3820: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 3821: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 3822: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3823: 	bneq	%r1, %r2, bneq_else.9017
"11001100000000010000000000000001",	-- 3824: 	lli	%r1, 1
"01010100000000000000111011110011",	-- 3825: 	j	bneq_cont.9018
	-- bneq_else.9017:
"11001100000000010000000000000000",	-- 3826: 	lli	%r1, 0
	-- bneq_cont.9018:
	-- bneq_cont.9016:
	-- bneq_cont.9014:
"11001100000000100000000000000000",	-- 3827: 	lli	%r2, 0
"00101000001000100000000001100011",	-- 3828: 	bneq	%r1, %r2, bneq_else.9019
"11001100000000010000000000000100",	-- 3829: 	lli	%r1, 4
"00111011110000100000000000000011",	-- 3830: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 3831: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3832: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000000100",	-- 3833: 	lf	%f1, [%sp + 4]
"11100100000000010000000000000000",	-- 3834: 	subf	%f0, %f0, %f1
"11001100000000010000000000000101",	-- 3835: 	lli	%r1, 5
"10000100010000010000100000000000",	-- 3836: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 3837: 	lf	%f1, [%r1 + 0]
"11101000000000010000000000000000",	-- 3838: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000000",	-- 3839: 	lli	%r1, 0
"00111011110000110000000000000110",	-- 3840: 	lw	%r3, [%sp + 6]
"10000100011000010000100000000000",	-- 3841: 	add	%r1, %r3, %r1
"10010000001000010000000000000000",	-- 3842: 	lf	%f1, [%r1 + 0]
"11101000000000010000100000000000",	-- 3843: 	mulf	%f1, %f0, %f1
"10010011110000100000000000000001",	-- 3844: 	lf	%f2, [%sp + 1]
"11100000001000100000100000000000",	-- 3845: 	addf	%f1, %f1, %f2
"10110000000111100000000000001101",	-- 3846: 	sf	%f0, [%sp + 13]
"00001100001000000000000000000000",	-- 3847: 	movf	%f0, %f1
"00111111111111100000000000001110",	-- 3848: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 3849: 	addi	%sp, %sp, 15
"01011000000000000010101001001111",	-- 3850: 	jal	yj_fabs
"10101011110111100000000000001111",	-- 3851: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 3852: 	lw	%ra, [%sp + 14]
"00111011110000010000000000000111",	-- 3853: 	lw	%r1, [%sp + 7]
"10110000000111100000000000001110",	-- 3854: 	sf	%f0, [%sp + 14]
"00111111111111100000000000001111",	-- 3855: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 3856: 	addi	%sp, %sp, 16
"01011000000000000000011001011010",	-- 3857: 	jal	o_param_a.2632
"10101011110111100000000000010000",	-- 3858: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 3859: 	lw	%ra, [%sp + 15]
"00001100000000010000000000000000",	-- 3860: 	movf	%f1, %f0
"10010011110000000000000000001110",	-- 3861: 	lf	%f0, [%sp + 14]
"00111111111111100000000000001111",	-- 3862: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 3863: 	addi	%sp, %sp, 16
"01011000000000000000010011110011",	-- 3864: 	jal	fless.2532
"10101011110111100000000000010000",	-- 3865: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 3866: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 3867: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3868: 	bneq	%r1, %r2, bneq_else.9020
"11001100000000010000000000000000",	-- 3869: 	lli	%r1, 0
"01010100000000000000111101001100",	-- 3870: 	j	bneq_cont.9021
	-- bneq_else.9020:
"11001100000000010000000000000001",	-- 3871: 	lli	%r1, 1
"00111011110000100000000000000110",	-- 3872: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 3873: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3874: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000001101",	-- 3875: 	lf	%f1, [%sp + 13]
"11101000001000000000000000000000",	-- 3876: 	mulf	%f0, %f1, %f0
"10010011110000100000000000000010",	-- 3877: 	lf	%f2, [%sp + 2]
"11100000000000100000000000000000",	-- 3878: 	addf	%f0, %f0, %f2
"00111111111111100000000000001111",	-- 3879: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 3880: 	addi	%sp, %sp, 16
"01011000000000000010101001001111",	-- 3881: 	jal	yj_fabs
"10101011110111100000000000010000",	-- 3882: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 3883: 	lw	%ra, [%sp + 15]
"00111011110000010000000000000111",	-- 3884: 	lw	%r1, [%sp + 7]
"10110000000111100000000000001111",	-- 3885: 	sf	%f0, [%sp + 15]
"00111111111111100000000000010000",	-- 3886: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 3887: 	addi	%sp, %sp, 17
"01011000000000000000011001011111",	-- 3888: 	jal	o_param_b.2634
"10101011110111100000000000010001",	-- 3889: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 3890: 	lw	%ra, [%sp + 16]
"00001100000000010000000000000000",	-- 3891: 	movf	%f1, %f0
"10010011110000000000000000001111",	-- 3892: 	lf	%f0, [%sp + 15]
"00111111111111100000000000010000",	-- 3893: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 3894: 	addi	%sp, %sp, 17
"01011000000000000000010011110011",	-- 3895: 	jal	fless.2532
"10101011110111100000000000010001",	-- 3896: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 3897: 	lw	%ra, [%sp + 16]
"11001100000000100000000000000000",	-- 3898: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3899: 	bneq	%r1, %r2, bneq_else.9022
"11001100000000010000000000000000",	-- 3900: 	lli	%r1, 0
"01010100000000000000111101001100",	-- 3901: 	j	bneq_cont.9023
	-- bneq_else.9022:
"11001100000000010000000000000101",	-- 3902: 	lli	%r1, 5
"00111011110000100000000000000011",	-- 3903: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 3904: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 3905: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000010000",	-- 3906: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 3907: 	addi	%sp, %sp, 17
"01011000000000000000010011100100",	-- 3908: 	jal	fiszero.2526
"10101011110111100000000000010001",	-- 3909: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 3910: 	lw	%ra, [%sp + 16]
"11001100000000100000000000000000",	-- 3911: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3912: 	bneq	%r1, %r2, bneq_else.9024
"11001100000000010000000000000001",	-- 3913: 	lli	%r1, 1
"01010100000000000000111101001100",	-- 3914: 	j	bneq_cont.9025
	-- bneq_else.9024:
"11001100000000010000000000000000",	-- 3915: 	lli	%r1, 0
	-- bneq_cont.9025:
	-- bneq_cont.9023:
	-- bneq_cont.9021:
"11001100000000100000000000000000",	-- 3916: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3917: 	bneq	%r1, %r2, bneq_else.9026
"11001100000000010000000000000000",	-- 3918: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3919: 	jr	%ra
	-- bneq_else.9026:
"11001100000000010000000000000000",	-- 3920: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 3921: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3922: 	add	%r1, %r2, %r1
"10010011110000000000000000001101",	-- 3923: 	lf	%f0, [%sp + 13]
"10110000000000010000000000000000",	-- 3924: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 3925: 	lli	%r1, 3
"01001111111000000000000000000000",	-- 3926: 	jr	%ra
	-- bneq_else.9019:
"11001100000000010000000000000000",	-- 3927: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 3928: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3929: 	add	%r1, %r2, %r1
"10010011110000000000000000001010",	-- 3930: 	lf	%f0, [%sp + 10]
"10110000000000010000000000000000",	-- 3931: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 3932: 	lli	%r1, 2
"01001111111000000000000000000000",	-- 3933: 	jr	%ra
	-- bneq_else.9012:
"11001100000000010000000000000000",	-- 3934: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 3935: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3936: 	add	%r1, %r2, %r1
"10010011110000000000000000000101",	-- 3937: 	lf	%f0, [%sp + 5]
"10110000000000010000000000000000",	-- 3938: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 3939: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 3940: 	jr	%ra
	-- solver_surface_fast.2767:
"00111011011000010000000000000001",	-- 3941: 	lw	%r1, [%r27 + 1]
"11001100000000110000000000000000",	-- 3942: 	lli	%r3, 0
"10000100010000110001100000000000",	-- 3943: 	add	%r3, %r2, %r3
"10010000011000110000000000000000",	-- 3944: 	lf	%f3, [%r3 + 0]
"00111100001111100000000000000000",	-- 3945: 	sw	%r1, [%sp + 0]
"10110000010111100000000000000001",	-- 3946: 	sf	%f2, [%sp + 1]
"10110000001111100000000000000010",	-- 3947: 	sf	%f1, [%sp + 2]
"10110000000111100000000000000011",	-- 3948: 	sf	%f0, [%sp + 3]
"00111100010111100000000000000100",	-- 3949: 	sw	%r2, [%sp + 4]
"00001100011000000000000000000000",	-- 3950: 	movf	%f0, %f3
"00111111111111100000000000000101",	-- 3951: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 3952: 	addi	%sp, %sp, 6
"01011000000000000000010011011101",	-- 3953: 	jal	fisneg.2524
"10101011110111100000000000000110",	-- 3954: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 3955: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000000",	-- 3956: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 3957: 	bneq	%r1, %r2, bneq_else.9027
"11001100000000010000000000000000",	-- 3958: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 3959: 	jr	%ra
	-- bneq_else.9027:
"11001100000000010000000000000000",	-- 3960: 	lli	%r1, 0
"11001100000000100000000000000001",	-- 3961: 	lli	%r2, 1
"00111011110000110000000000000100",	-- 3962: 	lw	%r3, [%sp + 4]
"10000100011000100001000000000000",	-- 3963: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 3964: 	lf	%f0, [%r2 + 0]
"10010011110000010000000000000011",	-- 3965: 	lf	%f1, [%sp + 3]
"11101000000000010000000000000000",	-- 3966: 	mulf	%f0, %f0, %f1
"11001100000000100000000000000010",	-- 3967: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 3968: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 3969: 	lf	%f1, [%r2 + 0]
"10010011110000100000000000000010",	-- 3970: 	lf	%f2, [%sp + 2]
"11101000001000100000100000000000",	-- 3971: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 3972: 	addf	%f0, %f0, %f1
"11001100000000100000000000000011",	-- 3973: 	lli	%r2, 3
"10000100011000100001000000000000",	-- 3974: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 3975: 	lf	%f1, [%r2 + 0]
"10010011110000100000000000000001",	-- 3976: 	lf	%f2, [%sp + 1]
"11101000001000100000100000000000",	-- 3977: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 3978: 	addf	%f0, %f0, %f1
"00111011110000100000000000000000",	-- 3979: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 3980: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 3981: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 3982: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 3983: 	jr	%ra
	-- solver_second_fast.2773:
"00111011011000110000000000000001",	-- 3984: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 3985: 	lli	%r4, 0
"10000100010001000010000000000000",	-- 3986: 	add	%r4, %r2, %r4
"10010000100000110000000000000000",	-- 3987: 	lf	%f3, [%r4 + 0]
"00111100011111100000000000000000",	-- 3988: 	sw	%r3, [%sp + 0]
"10110000011111100000000000000001",	-- 3989: 	sf	%f3, [%sp + 1]
"00111100001111100000000000000010",	-- 3990: 	sw	%r1, [%sp + 2]
"10110000010111100000000000000011",	-- 3991: 	sf	%f2, [%sp + 3]
"10110000001111100000000000000100",	-- 3992: 	sf	%f1, [%sp + 4]
"10110000000111100000000000000101",	-- 3993: 	sf	%f0, [%sp + 5]
"00111100010111100000000000000110",	-- 3994: 	sw	%r2, [%sp + 6]
"00001100011000000000000000000000",	-- 3995: 	movf	%f0, %f3
"00111111111111100000000000000111",	-- 3996: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 3997: 	addi	%sp, %sp, 8
"01011000000000000000010011100100",	-- 3998: 	jal	fiszero.2526
"10101011110111100000000000001000",	-- 3999: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 4000: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000000",	-- 4001: 	lli	%r2, 0
"00101000001000100000000001110011",	-- 4002: 	bneq	%r1, %r2, bneq_else.9028
"11001100000000010000000000000001",	-- 4003: 	lli	%r1, 1
"00111011110000100000000000000110",	-- 4004: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 4005: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 4006: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000000101",	-- 4007: 	lf	%f1, [%sp + 5]
"11101000000000010000000000000000",	-- 4008: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000010",	-- 4009: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 4010: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 4011: 	lf	%f2, [%r1 + 0]
"10010011110000110000000000000100",	-- 4012: 	lf	%f3, [%sp + 4]
"11101000010000110001000000000000",	-- 4013: 	mulf	%f2, %f2, %f3
"11100000000000100000000000000000",	-- 4014: 	addf	%f0, %f0, %f2
"11001100000000010000000000000011",	-- 4015: 	lli	%r1, 3
"10000100010000010000100000000000",	-- 4016: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 4017: 	lf	%f2, [%r1 + 0]
"10010011110001000000000000000011",	-- 4018: 	lf	%f4, [%sp + 3]
"11101000010001000001000000000000",	-- 4019: 	mulf	%f2, %f2, %f4
"11100000000000100000000000000000",	-- 4020: 	addf	%f0, %f0, %f2
"00111011110000010000000000000010",	-- 4021: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000111",	-- 4022: 	sf	%f0, [%sp + 7]
"00001100100000100000000000000000",	-- 4023: 	movf	%f2, %f4
"00001100001000000000000000000000",	-- 4024: 	movf	%f0, %f1
"00001100011000010000000000000000",	-- 4025: 	movf	%f1, %f3
"00111111111111100000000000001000",	-- 4026: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 4027: 	addi	%sp, %sp, 9
"01011000000000000000110001111010",	-- 4028: 	jal	quadratic.2737
"10101011110111100000000000001001",	-- 4029: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 4030: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000010",	-- 4031: 	lw	%r1, [%sp + 2]
"10110000000111100000000000001000",	-- 4032: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 4033: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4034: 	addi	%sp, %sp, 10
"01011000000000000000011001010010",	-- 4035: 	jal	o_form.2624
"10101011110111100000000000001010",	-- 4036: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4037: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000011",	-- 4038: 	lli	%r2, 3
"00101000001000100000000000000110",	-- 4039: 	bneq	%r1, %r2, bneq_else.9029
"00010100000000000000000000000000",	-- 4040: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 4041: 	lhif	%f0, 1.000000
"10010011110000010000000000001000",	-- 4042: 	lf	%f1, [%sp + 8]
"11100100001000000000000000000000",	-- 4043: 	subf	%f0, %f1, %f0
"01010100000000000000111111001110",	-- 4044: 	j	bneq_cont.9030
	-- bneq_else.9029:
"10010011110000000000000000001000",	-- 4045: 	lf	%f0, [%sp + 8]
	-- bneq_cont.9030:
"10010011110000010000000000000111",	-- 4046: 	lf	%f1, [%sp + 7]
"10110000000111100000000000001001",	-- 4047: 	sf	%f0, [%sp + 9]
"00001100001000000000000000000000",	-- 4048: 	movf	%f0, %f1
"00111111111111100000000000001010",	-- 4049: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4050: 	addi	%sp, %sp, 11
"01011000000000000000010011110001",	-- 4051: 	jal	fsqr.2530
"10101011110111100000000000001011",	-- 4052: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4053: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 4054: 	lf	%f1, [%sp + 9]
"10010011110000100000000000000001",	-- 4055: 	lf	%f2, [%sp + 1]
"11101000010000010000100000000000",	-- 4056: 	mulf	%f1, %f2, %f1
"11100100000000010000000000000000",	-- 4057: 	subf	%f0, %f0, %f1
"10110000000111100000000000001010",	-- 4058: 	sf	%f0, [%sp + 10]
"00111111111111100000000000001011",	-- 4059: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4060: 	addi	%sp, %sp, 12
"01011000000000000000010011010110",	-- 4061: 	jal	fispos.2522
"10101011110111100000000000001100",	-- 4062: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4063: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 4064: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 4065: 	bneq	%r1, %r2, bneq_else.9031
"11001100000000010000000000000000",	-- 4066: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 4067: 	jr	%ra
	-- bneq_else.9031:
"00111011110000010000000000000010",	-- 4068: 	lw	%r1, [%sp + 2]
"00111111111111100000000000001011",	-- 4069: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4070: 	addi	%sp, %sp, 12
"01011000000000000000011001010110",	-- 4071: 	jal	o_isinvert.2628
"10101011110111100000000000001100",	-- 4072: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4073: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 4074: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 4075: 	bneq	%r1, %r2, bneq_else.9032
"11001100000000010000000000000000",	-- 4076: 	lli	%r1, 0
"10010011110000000000000000001010",	-- 4077: 	lf	%f0, [%sp + 10]
"00111100001111100000000000001011",	-- 4078: 	sw	%r1, [%sp + 11]
"00111111111111100000000000001100",	-- 4079: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4080: 	addi	%sp, %sp, 13
"01011000000000000010101000110000",	-- 4081: 	jal	yj_sqrt
"10101011110111100000000000001101",	-- 4082: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4083: 	lw	%ra, [%sp + 12]
"10010011110000010000000000000111",	-- 4084: 	lf	%f1, [%sp + 7]
"11100100001000000000000000000000",	-- 4085: 	subf	%f0, %f1, %f0
"11001100000000010000000000000100",	-- 4086: 	lli	%r1, 4
"00111011110000100000000000000110",	-- 4087: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 4088: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4089: 	lf	%f1, [%r1 + 0]
"11101000000000010000000000000000",	-- 4090: 	mulf	%f0, %f0, %f1
"00111011110000010000000000001011",	-- 4091: 	lw	%r1, [%sp + 11]
"00111011110000100000000000000000",	-- 4092: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 4093: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4094: 	sf	%f0, [%r1 + 0]
"01010100000000000001000000010011",	-- 4095: 	j	bneq_cont.9033
	-- bneq_else.9032:
"11001100000000010000000000000000",	-- 4096: 	lli	%r1, 0
"10010011110000000000000000001010",	-- 4097: 	lf	%f0, [%sp + 10]
"00111100001111100000000000001100",	-- 4098: 	sw	%r1, [%sp + 12]
"00111111111111100000000000001101",	-- 4099: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 4100: 	addi	%sp, %sp, 14
"01011000000000000010101000110000",	-- 4101: 	jal	yj_sqrt
"10101011110111100000000000001110",	-- 4102: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 4103: 	lw	%ra, [%sp + 13]
"10010011110000010000000000000111",	-- 4104: 	lf	%f1, [%sp + 7]
"11100000001000000000000000000000",	-- 4105: 	addf	%f0, %f1, %f0
"11001100000000010000000000000100",	-- 4106: 	lli	%r1, 4
"00111011110000100000000000000110",	-- 4107: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 4108: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4109: 	lf	%f1, [%r1 + 0]
"11101000000000010000000000000000",	-- 4110: 	mulf	%f0, %f0, %f1
"00111011110000010000000000001100",	-- 4111: 	lw	%r1, [%sp + 12]
"00111011110000100000000000000000",	-- 4112: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 4113: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4114: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9033:
"11001100000000010000000000000001",	-- 4115: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 4116: 	jr	%ra
	-- bneq_else.9028:
"11001100000000010000000000000000",	-- 4117: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 4118: 	jr	%ra
	-- solver_fast.2779:
"00111011011001000000000000000100",	-- 4119: 	lw	%r4, [%r27 + 4]
"00111011011001010000000000000011",	-- 4120: 	lw	%r5, [%r27 + 3]
"00111011011001100000000000000010",	-- 4121: 	lw	%r6, [%r27 + 2]
"00111011011001110000000000000001",	-- 4122: 	lw	%r7, [%r27 + 1]
"10000100111000010011100000000000",	-- 4123: 	add	%r7, %r7, %r1
"00111000111001110000000000000000",	-- 4124: 	lw	%r7, [%r7 + 0]
"11001100000010000000000000000000",	-- 4125: 	lli	%r8, 0
"10000100011010000100000000000000",	-- 4126: 	add	%r8, %r3, %r8
"10010001000000000000000000000000",	-- 4127: 	lf	%f0, [%r8 + 0]
"00111100101111100000000000000000",	-- 4128: 	sw	%r5, [%sp + 0]
"00111100100111100000000000000001",	-- 4129: 	sw	%r4, [%sp + 1]
"00111100110111100000000000000010",	-- 4130: 	sw	%r6, [%sp + 2]
"00111100001111100000000000000011",	-- 4131: 	sw	%r1, [%sp + 3]
"00111100010111100000000000000100",	-- 4132: 	sw	%r2, [%sp + 4]
"00111100111111100000000000000101",	-- 4133: 	sw	%r7, [%sp + 5]
"00111100011111100000000000000110",	-- 4134: 	sw	%r3, [%sp + 6]
"10110000000111100000000000000111",	-- 4135: 	sf	%f0, [%sp + 7]
"10000100000001110000100000000000",	-- 4136: 	add	%r1, %r0, %r7
"00111111111111100000000000001000",	-- 4137: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 4138: 	addi	%sp, %sp, 9
"01011000000000000000011001101011",	-- 4139: 	jal	o_param_x.2640
"10101011110111100000000000001001",	-- 4140: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 4141: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000111",	-- 4142: 	lf	%f1, [%sp + 7]
"11100100001000000000000000000000",	-- 4143: 	subf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 4144: 	lli	%r1, 1
"00111011110000100000000000000110",	-- 4145: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 4146: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4147: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000101",	-- 4148: 	lw	%r1, [%sp + 5]
"10110000000111100000000000001000",	-- 4149: 	sf	%f0, [%sp + 8]
"10110000001111100000000000001001",	-- 4150: 	sf	%f1, [%sp + 9]
"00111111111111100000000000001010",	-- 4151: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4152: 	addi	%sp, %sp, 11
"01011000000000000000011001110000",	-- 4153: 	jal	o_param_y.2642
"10101011110111100000000000001011",	-- 4154: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4155: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 4156: 	lf	%f1, [%sp + 9]
"11100100001000000000000000000000",	-- 4157: 	subf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 4158: 	lli	%r1, 2
"00111011110000100000000000000110",	-- 4159: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 4160: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4161: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000101",	-- 4162: 	lw	%r1, [%sp + 5]
"10110000000111100000000000001010",	-- 4163: 	sf	%f0, [%sp + 10]
"10110000001111100000000000001011",	-- 4164: 	sf	%f1, [%sp + 11]
"00111111111111100000000000001100",	-- 4165: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4166: 	addi	%sp, %sp, 13
"01011000000000000000011001110101",	-- 4167: 	jal	o_param_z.2644
"10101011110111100000000000001101",	-- 4168: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4169: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001011",	-- 4170: 	lf	%f1, [%sp + 11]
"11100100001000000000000000000000",	-- 4171: 	subf	%f0, %f1, %f0
"00111011110000010000000000000100",	-- 4172: 	lw	%r1, [%sp + 4]
"10110000000111100000000000001100",	-- 4173: 	sf	%f0, [%sp + 12]
"00111111111111100000000000001101",	-- 4174: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 4175: 	addi	%sp, %sp, 14
"01011000000000000000011010111110",	-- 4176: 	jal	d_const.2685
"10101011110111100000000000001110",	-- 4177: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 4178: 	lw	%ra, [%sp + 13]
"00111011110000100000000000000011",	-- 4179: 	lw	%r2, [%sp + 3]
"10000100001000100000100000000000",	-- 4180: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 4181: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000000101",	-- 4182: 	lw	%r2, [%sp + 5]
"00111100001111100000000000001101",	-- 4183: 	sw	%r1, [%sp + 13]
"10000100000000100000100000000000",	-- 4184: 	add	%r1, %r0, %r2
"00111111111111100000000000001110",	-- 4185: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 4186: 	addi	%sp, %sp, 15
"01011000000000000000011001010010",	-- 4187: 	jal	o_form.2624
"10101011110111100000000000001111",	-- 4188: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 4189: 	lw	%ra, [%sp + 14]
"11001100000000100000000000000001",	-- 4190: 	lli	%r2, 1
"00101000001000100000000000010000",	-- 4191: 	bneq	%r1, %r2, bneq_else.9034
"00111011110000010000000000000100",	-- 4192: 	lw	%r1, [%sp + 4]
"00111111111111100000000000001110",	-- 4193: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 4194: 	addi	%sp, %sp, 15
"01011000000000000000011010111100",	-- 4195: 	jal	d_vec.2683
"10101011110111100000000000001111",	-- 4196: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 4197: 	lw	%ra, [%sp + 14]
"10000100000000010001000000000000",	-- 4198: 	add	%r2, %r0, %r1
"10010011110000000000000000001000",	-- 4199: 	lf	%f0, [%sp + 8]
"10010011110000010000000000001010",	-- 4200: 	lf	%f1, [%sp + 10]
"10010011110000100000000000001100",	-- 4201: 	lf	%f2, [%sp + 12]
"00111011110000010000000000000101",	-- 4202: 	lw	%r1, [%sp + 5]
"00111011110000110000000000001101",	-- 4203: 	lw	%r3, [%sp + 13]
"00111011110110110000000000000010",	-- 4204: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 4205: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 4206: 	jr	%r26
	-- bneq_else.9034:
"11001100000000100000000000000010",	-- 4207: 	lli	%r2, 2
"00101000001000100000000000001001",	-- 4208: 	bneq	%r1, %r2, bneq_else.9035
"10010011110000000000000000001000",	-- 4209: 	lf	%f0, [%sp + 8]
"10010011110000010000000000001010",	-- 4210: 	lf	%f1, [%sp + 10]
"10010011110000100000000000001100",	-- 4211: 	lf	%f2, [%sp + 12]
"00111011110000010000000000000101",	-- 4212: 	lw	%r1, [%sp + 5]
"00111011110000100000000000001101",	-- 4213: 	lw	%r2, [%sp + 13]
"00111011110110110000000000000001",	-- 4214: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 4215: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 4216: 	jr	%r26
	-- bneq_else.9035:
"10010011110000000000000000001000",	-- 4217: 	lf	%f0, [%sp + 8]
"10010011110000010000000000001010",	-- 4218: 	lf	%f1, [%sp + 10]
"10010011110000100000000000001100",	-- 4219: 	lf	%f2, [%sp + 12]
"00111011110000010000000000000101",	-- 4220: 	lw	%r1, [%sp + 5]
"00111011110000100000000000001101",	-- 4221: 	lw	%r2, [%sp + 13]
"00111011110110110000000000000000",	-- 4222: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 4223: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 4224: 	jr	%r26
	-- solver_surface_fast2.2783:
"00111011011000010000000000000001",	-- 4225: 	lw	%r1, [%r27 + 1]
"11001100000001000000000000000000",	-- 4226: 	lli	%r4, 0
"10000100010001000010000000000000",	-- 4227: 	add	%r4, %r2, %r4
"10010000100000000000000000000000",	-- 4228: 	lf	%f0, [%r4 + 0]
"00111100001111100000000000000000",	-- 4229: 	sw	%r1, [%sp + 0]
"00111100011111100000000000000001",	-- 4230: 	sw	%r3, [%sp + 1]
"00111100010111100000000000000010",	-- 4231: 	sw	%r2, [%sp + 2]
"00111111111111100000000000000011",	-- 4232: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 4233: 	addi	%sp, %sp, 4
"01011000000000000000010011011101",	-- 4234: 	jal	fisneg.2524
"10101011110111100000000000000100",	-- 4235: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 4236: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000000",	-- 4237: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 4238: 	bneq	%r1, %r2, bneq_else.9036
"11001100000000010000000000000000",	-- 4239: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 4240: 	jr	%ra
	-- bneq_else.9036:
"11001100000000010000000000000000",	-- 4241: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 4242: 	lli	%r2, 0
"00111011110000110000000000000010",	-- 4243: 	lw	%r3, [%sp + 2]
"10000100011000100001000000000000",	-- 4244: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4245: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000011",	-- 4246: 	lli	%r2, 3
"00111011110000110000000000000001",	-- 4247: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4248: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 4249: 	lf	%f1, [%r2 + 0]
"11101000000000010000000000000000",	-- 4250: 	mulf	%f0, %f0, %f1
"00111011110000100000000000000000",	-- 4251: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 4252: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4253: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 4254: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 4255: 	jr	%ra
	-- solver_second_fast2.2790:
"00111011011001000000000000000001",	-- 4256: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 4257: 	lli	%r5, 0
"10000100010001010010100000000000",	-- 4258: 	add	%r5, %r2, %r5
"10010000101000110000000000000000",	-- 4259: 	lf	%f3, [%r5 + 0]
"00111100100111100000000000000000",	-- 4260: 	sw	%r4, [%sp + 0]
"00111100001111100000000000000001",	-- 4261: 	sw	%r1, [%sp + 1]
"10110000011111100000000000000010",	-- 4262: 	sf	%f3, [%sp + 2]
"00111100011111100000000000000011",	-- 4263: 	sw	%r3, [%sp + 3]
"10110000010111100000000000000100",	-- 4264: 	sf	%f2, [%sp + 4]
"10110000001111100000000000000101",	-- 4265: 	sf	%f1, [%sp + 5]
"10110000000111100000000000000110",	-- 4266: 	sf	%f0, [%sp + 6]
"00111100010111100000000000000111",	-- 4267: 	sw	%r2, [%sp + 7]
"00001100011000000000000000000000",	-- 4268: 	movf	%f0, %f3
"00111111111111100000000000001000",	-- 4269: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 4270: 	addi	%sp, %sp, 9
"01011000000000000000010011100100",	-- 4271: 	jal	fiszero.2526
"10101011110111100000000000001001",	-- 4272: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 4273: 	lw	%ra, [%sp + 8]
"11001100000000100000000000000000",	-- 4274: 	lli	%r2, 0
"00101000001000100000000001011101",	-- 4275: 	bneq	%r1, %r2, bneq_else.9037
"11001100000000010000000000000001",	-- 4276: 	lli	%r1, 1
"00111011110000100000000000000111",	-- 4277: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 4278: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 4279: 	lf	%f0, [%r1 + 0]
"10010011110000010000000000000110",	-- 4280: 	lf	%f1, [%sp + 6]
"11101000000000010000000000000000",	-- 4281: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000010",	-- 4282: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 4283: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4284: 	lf	%f1, [%r1 + 0]
"10010011110000100000000000000101",	-- 4285: 	lf	%f2, [%sp + 5]
"11101000001000100000100000000000",	-- 4286: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 4287: 	addf	%f0, %f0, %f1
"11001100000000010000000000000011",	-- 4288: 	lli	%r1, 3
"10000100010000010000100000000000",	-- 4289: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4290: 	lf	%f1, [%r1 + 0]
"10010011110000100000000000000100",	-- 4291: 	lf	%f2, [%sp + 4]
"11101000001000100000100000000000",	-- 4292: 	mulf	%f1, %f1, %f2
"11100000000000010000000000000000",	-- 4293: 	addf	%f0, %f0, %f1
"11001100000000010000000000000011",	-- 4294: 	lli	%r1, 3
"00111011110000110000000000000011",	-- 4295: 	lw	%r3, [%sp + 3]
"10000100011000010000100000000000",	-- 4296: 	add	%r1, %r3, %r1
"10010000001000010000000000000000",	-- 4297: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000001000",	-- 4298: 	sf	%f0, [%sp + 8]
"10110000001111100000000000001001",	-- 4299: 	sf	%f1, [%sp + 9]
"00111111111111100000000000001010",	-- 4300: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4301: 	addi	%sp, %sp, 11
"01011000000000000000010011110001",	-- 4302: 	jal	fsqr.2530
"10101011110111100000000000001011",	-- 4303: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4304: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 4305: 	lf	%f1, [%sp + 9]
"10010011110000100000000000000010",	-- 4306: 	lf	%f2, [%sp + 2]
"11101000010000010000100000000000",	-- 4307: 	mulf	%f1, %f2, %f1
"11100100000000010000000000000000",	-- 4308: 	subf	%f0, %f0, %f1
"10110000000111100000000000001010",	-- 4309: 	sf	%f0, [%sp + 10]
"00111111111111100000000000001011",	-- 4310: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4311: 	addi	%sp, %sp, 12
"01011000000000000000010011010110",	-- 4312: 	jal	fispos.2522
"10101011110111100000000000001100",	-- 4313: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4314: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 4315: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 4316: 	bneq	%r1, %r2, bneq_else.9038
"11001100000000010000000000000000",	-- 4317: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 4318: 	jr	%ra
	-- bneq_else.9038:
"00111011110000010000000000000001",	-- 4319: 	lw	%r1, [%sp + 1]
"00111111111111100000000000001011",	-- 4320: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4321: 	addi	%sp, %sp, 12
"01011000000000000000011001010110",	-- 4322: 	jal	o_isinvert.2628
"10101011110111100000000000001100",	-- 4323: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4324: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 4325: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 4326: 	bneq	%r1, %r2, bneq_else.9039
"11001100000000010000000000000000",	-- 4327: 	lli	%r1, 0
"10010011110000000000000000001010",	-- 4328: 	lf	%f0, [%sp + 10]
"00111100001111100000000000001011",	-- 4329: 	sw	%r1, [%sp + 11]
"00111111111111100000000000001100",	-- 4330: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4331: 	addi	%sp, %sp, 13
"01011000000000000010101000110000",	-- 4332: 	jal	yj_sqrt
"10101011110111100000000000001101",	-- 4333: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4334: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001000",	-- 4335: 	lf	%f1, [%sp + 8]
"11100100001000000000000000000000",	-- 4336: 	subf	%f0, %f1, %f0
"11001100000000010000000000000100",	-- 4337: 	lli	%r1, 4
"00111011110000100000000000000111",	-- 4338: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 4339: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4340: 	lf	%f1, [%r1 + 0]
"11101000000000010000000000000000",	-- 4341: 	mulf	%f0, %f0, %f1
"00111011110000010000000000001011",	-- 4342: 	lw	%r1, [%sp + 11]
"00111011110000100000000000000000",	-- 4343: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 4344: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4345: 	sf	%f0, [%r1 + 0]
"01010100000000000001000100001110",	-- 4346: 	j	bneq_cont.9040
	-- bneq_else.9039:
"11001100000000010000000000000000",	-- 4347: 	lli	%r1, 0
"10010011110000000000000000001010",	-- 4348: 	lf	%f0, [%sp + 10]
"00111100001111100000000000001100",	-- 4349: 	sw	%r1, [%sp + 12]
"00111111111111100000000000001101",	-- 4350: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 4351: 	addi	%sp, %sp, 14
"01011000000000000010101000110000",	-- 4352: 	jal	yj_sqrt
"10101011110111100000000000001110",	-- 4353: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 4354: 	lw	%ra, [%sp + 13]
"10010011110000010000000000001000",	-- 4355: 	lf	%f1, [%sp + 8]
"11100000001000000000000000000000",	-- 4356: 	addf	%f0, %f1, %f0
"11001100000000010000000000000100",	-- 4357: 	lli	%r1, 4
"00111011110000100000000000000111",	-- 4358: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 4359: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4360: 	lf	%f1, [%r1 + 0]
"11101000000000010000000000000000",	-- 4361: 	mulf	%f0, %f0, %f1
"00111011110000010000000000001100",	-- 4362: 	lw	%r1, [%sp + 12]
"00111011110000100000000000000000",	-- 4363: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 4364: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4365: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9040:
"11001100000000010000000000000001",	-- 4366: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 4367: 	jr	%ra
	-- bneq_else.9037:
"11001100000000010000000000000000",	-- 4368: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 4369: 	jr	%ra
	-- solver_fast2.2797:
"00111011011000110000000000000100",	-- 4370: 	lw	%r3, [%r27 + 4]
"00111011011001000000000000000011",	-- 4371: 	lw	%r4, [%r27 + 3]
"00111011011001010000000000000010",	-- 4372: 	lw	%r5, [%r27 + 2]
"00111011011001100000000000000001",	-- 4373: 	lw	%r6, [%r27 + 1]
"10000100110000010011000000000000",	-- 4374: 	add	%r6, %r6, %r1
"00111000110001100000000000000000",	-- 4375: 	lw	%r6, [%r6 + 0]
"00111100100111100000000000000000",	-- 4376: 	sw	%r4, [%sp + 0]
"00111100011111100000000000000001",	-- 4377: 	sw	%r3, [%sp + 1]
"00111100101111100000000000000010",	-- 4378: 	sw	%r5, [%sp + 2]
"00111100110111100000000000000011",	-- 4379: 	sw	%r6, [%sp + 3]
"00111100001111100000000000000100",	-- 4380: 	sw	%r1, [%sp + 4]
"00111100010111100000000000000101",	-- 4381: 	sw	%r2, [%sp + 5]
"10000100000001100000100000000000",	-- 4382: 	add	%r1, %r0, %r6
"00111111111111100000000000000110",	-- 4383: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 4384: 	addi	%sp, %sp, 7
"01011000000000000000011010100010",	-- 4385: 	jal	o_param_ctbl.2662
"10101011110111100000000000000111",	-- 4386: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 4387: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 4388: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 4389: 	add	%r2, %r1, %r2
"10010000010000000000000000000000",	-- 4390: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000001",	-- 4391: 	lli	%r2, 1
"10000100001000100001000000000000",	-- 4392: 	add	%r2, %r1, %r2
"10010000010000010000000000000000",	-- 4393: 	lf	%f1, [%r2 + 0]
"11001100000000100000000000000010",	-- 4394: 	lli	%r2, 2
"10000100001000100001000000000000",	-- 4395: 	add	%r2, %r1, %r2
"10010000010000100000000000000000",	-- 4396: 	lf	%f2, [%r2 + 0]
"00111011110000100000000000000101",	-- 4397: 	lw	%r2, [%sp + 5]
"00111100001111100000000000000110",	-- 4398: 	sw	%r1, [%sp + 6]
"10110000010111100000000000000111",	-- 4399: 	sf	%f2, [%sp + 7]
"10110000001111100000000000001000",	-- 4400: 	sf	%f1, [%sp + 8]
"10110000000111100000000000001001",	-- 4401: 	sf	%f0, [%sp + 9]
"10000100000000100000100000000000",	-- 4402: 	add	%r1, %r0, %r2
"00111111111111100000000000001010",	-- 4403: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4404: 	addi	%sp, %sp, 11
"01011000000000000000011010111110",	-- 4405: 	jal	d_const.2685
"10101011110111100000000000001011",	-- 4406: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4407: 	lw	%ra, [%sp + 10]
"00111011110000100000000000000100",	-- 4408: 	lw	%r2, [%sp + 4]
"10000100001000100000100000000000",	-- 4409: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 4410: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000000011",	-- 4411: 	lw	%r2, [%sp + 3]
"00111100001111100000000000001010",	-- 4412: 	sw	%r1, [%sp + 10]
"10000100000000100000100000000000",	-- 4413: 	add	%r1, %r0, %r2
"00111111111111100000000000001011",	-- 4414: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4415: 	addi	%sp, %sp, 12
"01011000000000000000011001010010",	-- 4416: 	jal	o_form.2624
"10101011110111100000000000001100",	-- 4417: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4418: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000001",	-- 4419: 	lli	%r2, 1
"00101000001000100000000000010000",	-- 4420: 	bneq	%r1, %r2, bneq_else.9041
"00111011110000010000000000000101",	-- 4421: 	lw	%r1, [%sp + 5]
"00111111111111100000000000001011",	-- 4422: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4423: 	addi	%sp, %sp, 12
"01011000000000000000011010111100",	-- 4424: 	jal	d_vec.2683
"10101011110111100000000000001100",	-- 4425: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4426: 	lw	%ra, [%sp + 11]
"10000100000000010001000000000000",	-- 4427: 	add	%r2, %r0, %r1
"10010011110000000000000000001001",	-- 4428: 	lf	%f0, [%sp + 9]
"10010011110000010000000000001000",	-- 4429: 	lf	%f1, [%sp + 8]
"10010011110000100000000000000111",	-- 4430: 	lf	%f2, [%sp + 7]
"00111011110000010000000000000011",	-- 4431: 	lw	%r1, [%sp + 3]
"00111011110000110000000000001010",	-- 4432: 	lw	%r3, [%sp + 10]
"00111011110110110000000000000010",	-- 4433: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 4434: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 4435: 	jr	%r26
	-- bneq_else.9041:
"11001100000000100000000000000010",	-- 4436: 	lli	%r2, 2
"00101000001000100000000000001010",	-- 4437: 	bneq	%r1, %r2, bneq_else.9042
"10010011110000000000000000001001",	-- 4438: 	lf	%f0, [%sp + 9]
"10010011110000010000000000001000",	-- 4439: 	lf	%f1, [%sp + 8]
"10010011110000100000000000000111",	-- 4440: 	lf	%f2, [%sp + 7]
"00111011110000010000000000000011",	-- 4441: 	lw	%r1, [%sp + 3]
"00111011110000100000000000001010",	-- 4442: 	lw	%r2, [%sp + 10]
"00111011110000110000000000000110",	-- 4443: 	lw	%r3, [%sp + 6]
"00111011110110110000000000000001",	-- 4444: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 4445: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 4446: 	jr	%r26
	-- bneq_else.9042:
"10010011110000000000000000001001",	-- 4447: 	lf	%f0, [%sp + 9]
"10010011110000010000000000001000",	-- 4448: 	lf	%f1, [%sp + 8]
"10010011110000100000000000000111",	-- 4449: 	lf	%f2, [%sp + 7]
"00111011110000010000000000000011",	-- 4450: 	lw	%r1, [%sp + 3]
"00111011110000100000000000001010",	-- 4451: 	lw	%r2, [%sp + 10]
"00111011110000110000000000000110",	-- 4452: 	lw	%r3, [%sp + 6]
"00111011110110110000000000000000",	-- 4453: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 4454: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 4455: 	jr	%r26
	-- setup_rect_table.2800:
"11001100000000110000000000000110",	-- 4456: 	lli	%r3, 6
"00010100000000000000000000000000",	-- 4457: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4458: 	lhif	%f0, 0.000000
"00111100010111100000000000000000",	-- 4459: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 4460: 	sw	%r1, [%sp + 1]
"10000100000000110000100000000000",	-- 4461: 	add	%r1, %r0, %r3
"00111111111111100000000000000010",	-- 4462: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 4463: 	addi	%sp, %sp, 3
"01011000000000000010101000100100",	-- 4464: 	jal	yj_create_float_array
"10101011110111100000000000000011",	-- 4465: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 4466: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000000",	-- 4467: 	lli	%r2, 0
"00111011110000110000000000000001",	-- 4468: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4469: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4470: 	lf	%f0, [%r2 + 0]
"00111100001111100000000000000010",	-- 4471: 	sw	%r1, [%sp + 2]
"00111111111111100000000000000011",	-- 4472: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 4473: 	addi	%sp, %sp, 4
"01011000000000000000010011100100",	-- 4474: 	jal	fiszero.2526
"10101011110111100000000000000100",	-- 4475: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 4476: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000000",	-- 4477: 	lli	%r2, 0
"00101000001000100000000000111000",	-- 4478: 	bneq	%r1, %r2, bneq_else.9043
"11001100000000010000000000000000",	-- 4479: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 4480: 	lw	%r2, [%sp + 0]
"00111100001111100000000000000011",	-- 4481: 	sw	%r1, [%sp + 3]
"10000100000000100000100000000000",	-- 4482: 	add	%r1, %r0, %r2
"00111111111111100000000000000100",	-- 4483: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 4484: 	addi	%sp, %sp, 5
"01011000000000000000011001010110",	-- 4485: 	jal	o_isinvert.2628
"10101011110111100000000000000101",	-- 4486: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 4487: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000000",	-- 4488: 	lli	%r2, 0
"00111011110000110000000000000001",	-- 4489: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4490: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4491: 	lf	%f0, [%r2 + 0]
"00111100001111100000000000000100",	-- 4492: 	sw	%r1, [%sp + 4]
"00111111111111100000000000000101",	-- 4493: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 4494: 	addi	%sp, %sp, 6
"01011000000000000000010011011101",	-- 4495: 	jal	fisneg.2524
"10101011110111100000000000000110",	-- 4496: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 4497: 	lw	%ra, [%sp + 5]
"10000100000000010001000000000000",	-- 4498: 	add	%r2, %r0, %r1
"00111011110000010000000000000100",	-- 4499: 	lw	%r1, [%sp + 4]
"00111111111111100000000000000101",	-- 4500: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 4501: 	addi	%sp, %sp, 6
"01011000000000000000010011111000",	-- 4502: 	jal	xor.2565
"10101011110111100000000000000110",	-- 4503: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 4504: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000000",	-- 4505: 	lw	%r2, [%sp + 0]
"00111100001111100000000000000101",	-- 4506: 	sw	%r1, [%sp + 5]
"10000100000000100000100000000000",	-- 4507: 	add	%r1, %r0, %r2
"00111111111111100000000000000110",	-- 4508: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 4509: 	addi	%sp, %sp, 7
"01011000000000000000011001011010",	-- 4510: 	jal	o_param_a.2632
"10101011110111100000000000000111",	-- 4511: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 4512: 	lw	%ra, [%sp + 6]
"00111011110000010000000000000101",	-- 4513: 	lw	%r1, [%sp + 5]
"00111111111111100000000000000110",	-- 4514: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 4515: 	addi	%sp, %sp, 7
"01011000000000000000010100011011",	-- 4516: 	jal	fneg_cond.2570
"10101011110111100000000000000111",	-- 4517: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 4518: 	lw	%ra, [%sp + 6]
"00111011110000010000000000000011",	-- 4519: 	lw	%r1, [%sp + 3]
"00111011110000100000000000000010",	-- 4520: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4521: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4522: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 4523: 	lli	%r1, 1
"00010100000000000000000000000000",	-- 4524: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 4525: 	lhif	%f0, 1.000000
"11001100000000110000000000000000",	-- 4526: 	lli	%r3, 0
"00111011110001000000000000000001",	-- 4527: 	lw	%r4, [%sp + 1]
"10000100100000110001100000000000",	-- 4528: 	add	%r3, %r4, %r3
"10010000011000010000000000000000",	-- 4529: 	lf	%f1, [%r3 + 0]
"11101100000000010000000000000000",	-- 4530: 	divf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 4531: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4532: 	sf	%f0, [%r1 + 0]
"01010100000000000001000110111100",	-- 4533: 	j	bneq_cont.9044
	-- bneq_else.9043:
"11001100000000010000000000000001",	-- 4534: 	lli	%r1, 1
"00010100000000000000000000000000",	-- 4535: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4536: 	lhif	%f0, 0.000000
"00111011110000100000000000000010",	-- 4537: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4538: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4539: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9044:
"11001100000000010000000000000001",	-- 4540: 	lli	%r1, 1
"00111011110000110000000000000001",	-- 4541: 	lw	%r3, [%sp + 1]
"10000100011000010000100000000000",	-- 4542: 	add	%r1, %r3, %r1
"10010000001000000000000000000000",	-- 4543: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000000110",	-- 4544: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 4545: 	addi	%sp, %sp, 7
"01011000000000000000010011100100",	-- 4546: 	jal	fiszero.2526
"10101011110111100000000000000111",	-- 4547: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 4548: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 4549: 	lli	%r2, 0
"00101000001000100000000000111000",	-- 4550: 	bneq	%r1, %r2, bneq_else.9045
"11001100000000010000000000000010",	-- 4551: 	lli	%r1, 2
"00111011110000100000000000000000",	-- 4552: 	lw	%r2, [%sp + 0]
"00111100001111100000000000000110",	-- 4553: 	sw	%r1, [%sp + 6]
"10000100000000100000100000000000",	-- 4554: 	add	%r1, %r0, %r2
"00111111111111100000000000000111",	-- 4555: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 4556: 	addi	%sp, %sp, 8
"01011000000000000000011001010110",	-- 4557: 	jal	o_isinvert.2628
"10101011110111100000000000001000",	-- 4558: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 4559: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000001",	-- 4560: 	lli	%r2, 1
"00111011110000110000000000000001",	-- 4561: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4562: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4563: 	lf	%f0, [%r2 + 0]
"00111100001111100000000000000111",	-- 4564: 	sw	%r1, [%sp + 7]
"00111111111111100000000000001000",	-- 4565: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 4566: 	addi	%sp, %sp, 9
"01011000000000000000010011011101",	-- 4567: 	jal	fisneg.2524
"10101011110111100000000000001001",	-- 4568: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 4569: 	lw	%ra, [%sp + 8]
"10000100000000010001000000000000",	-- 4570: 	add	%r2, %r0, %r1
"00111011110000010000000000000111",	-- 4571: 	lw	%r1, [%sp + 7]
"00111111111111100000000000001000",	-- 4572: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 4573: 	addi	%sp, %sp, 9
"01011000000000000000010011111000",	-- 4574: 	jal	xor.2565
"10101011110111100000000000001001",	-- 4575: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 4576: 	lw	%ra, [%sp + 8]
"00111011110000100000000000000000",	-- 4577: 	lw	%r2, [%sp + 0]
"00111100001111100000000000001000",	-- 4578: 	sw	%r1, [%sp + 8]
"10000100000000100000100000000000",	-- 4579: 	add	%r1, %r0, %r2
"00111111111111100000000000001001",	-- 4580: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4581: 	addi	%sp, %sp, 10
"01011000000000000000011001011111",	-- 4582: 	jal	o_param_b.2634
"10101011110111100000000000001010",	-- 4583: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4584: 	lw	%ra, [%sp + 9]
"00111011110000010000000000001000",	-- 4585: 	lw	%r1, [%sp + 8]
"00111111111111100000000000001001",	-- 4586: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4587: 	addi	%sp, %sp, 10
"01011000000000000000010100011011",	-- 4588: 	jal	fneg_cond.2570
"10101011110111100000000000001010",	-- 4589: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4590: 	lw	%ra, [%sp + 9]
"00111011110000010000000000000110",	-- 4591: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000010",	-- 4592: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4593: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4594: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 4595: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 4596: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 4597: 	lhif	%f0, 1.000000
"11001100000000110000000000000001",	-- 4598: 	lli	%r3, 1
"00111011110001000000000000000001",	-- 4599: 	lw	%r4, [%sp + 1]
"10000100100000110001100000000000",	-- 4600: 	add	%r3, %r4, %r3
"10010000011000010000000000000000",	-- 4601: 	lf	%f1, [%r3 + 0]
"11101100000000010000000000000000",	-- 4602: 	divf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 4603: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4604: 	sf	%f0, [%r1 + 0]
"01010100000000000001001000000100",	-- 4605: 	j	bneq_cont.9046
	-- bneq_else.9045:
"11001100000000010000000000000011",	-- 4606: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 4607: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4608: 	lhif	%f0, 0.000000
"00111011110000100000000000000010",	-- 4609: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4610: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4611: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9046:
"11001100000000010000000000000010",	-- 4612: 	lli	%r1, 2
"00111011110000110000000000000001",	-- 4613: 	lw	%r3, [%sp + 1]
"10000100011000010000100000000000",	-- 4614: 	add	%r1, %r3, %r1
"10010000001000000000000000000000",	-- 4615: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000001001",	-- 4616: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4617: 	addi	%sp, %sp, 10
"01011000000000000000010011100100",	-- 4618: 	jal	fiszero.2526
"10101011110111100000000000001010",	-- 4619: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4620: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000000",	-- 4621: 	lli	%r2, 0
"00101000001000100000000000111000",	-- 4622: 	bneq	%r1, %r2, bneq_else.9047
"11001100000000010000000000000100",	-- 4623: 	lli	%r1, 4
"00111011110000100000000000000000",	-- 4624: 	lw	%r2, [%sp + 0]
"00111100001111100000000000001001",	-- 4625: 	sw	%r1, [%sp + 9]
"10000100000000100000100000000000",	-- 4626: 	add	%r1, %r0, %r2
"00111111111111100000000000001010",	-- 4627: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4628: 	addi	%sp, %sp, 11
"01011000000000000000011001010110",	-- 4629: 	jal	o_isinvert.2628
"10101011110111100000000000001011",	-- 4630: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4631: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000010",	-- 4632: 	lli	%r2, 2
"00111011110000110000000000000001",	-- 4633: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4634: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4635: 	lf	%f0, [%r2 + 0]
"00111100001111100000000000001010",	-- 4636: 	sw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 4637: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4638: 	addi	%sp, %sp, 12
"01011000000000000000010011011101",	-- 4639: 	jal	fisneg.2524
"10101011110111100000000000001100",	-- 4640: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4641: 	lw	%ra, [%sp + 11]
"10000100000000010001000000000000",	-- 4642: 	add	%r2, %r0, %r1
"00111011110000010000000000001010",	-- 4643: 	lw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 4644: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4645: 	addi	%sp, %sp, 12
"01011000000000000000010011111000",	-- 4646: 	jal	xor.2565
"10101011110111100000000000001100",	-- 4647: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4648: 	lw	%ra, [%sp + 11]
"00111011110000100000000000000000",	-- 4649: 	lw	%r2, [%sp + 0]
"00111100001111100000000000001011",	-- 4650: 	sw	%r1, [%sp + 11]
"10000100000000100000100000000000",	-- 4651: 	add	%r1, %r0, %r2
"00111111111111100000000000001100",	-- 4652: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4653: 	addi	%sp, %sp, 13
"01011000000000000000011001100100",	-- 4654: 	jal	o_param_c.2636
"10101011110111100000000000001101",	-- 4655: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4656: 	lw	%ra, [%sp + 12]
"00111011110000010000000000001011",	-- 4657: 	lw	%r1, [%sp + 11]
"00111111111111100000000000001100",	-- 4658: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4659: 	addi	%sp, %sp, 13
"01011000000000000000010100011011",	-- 4660: 	jal	fneg_cond.2570
"10101011110111100000000000001101",	-- 4661: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4662: 	lw	%ra, [%sp + 12]
"00111011110000010000000000001001",	-- 4663: 	lw	%r1, [%sp + 9]
"00111011110000100000000000000010",	-- 4664: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4665: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4666: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000101",	-- 4667: 	lli	%r1, 5
"00010100000000000000000000000000",	-- 4668: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 4669: 	lhif	%f0, 1.000000
"11001100000000110000000000000010",	-- 4670: 	lli	%r3, 2
"00111011110001000000000000000001",	-- 4671: 	lw	%r4, [%sp + 1]
"10000100100000110001100000000000",	-- 4672: 	add	%r3, %r4, %r3
"10010000011000010000000000000000",	-- 4673: 	lf	%f1, [%r3 + 0]
"11101100000000010000000000000000",	-- 4674: 	divf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 4675: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4676: 	sf	%f0, [%r1 + 0]
"01010100000000000001001001001100",	-- 4677: 	j	bneq_cont.9048
	-- bneq_else.9047:
"11001100000000010000000000000101",	-- 4678: 	lli	%r1, 5
"00010100000000000000000000000000",	-- 4679: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4680: 	lhif	%f0, 0.000000
"00111011110000100000000000000010",	-- 4681: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4682: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4683: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9048:
"10000100000000100000100000000000",	-- 4684: 	add	%r1, %r0, %r2
"01001111111000000000000000000000",	-- 4685: 	jr	%ra
	-- setup_surface_table.2803:
"11001100000000110000000000000100",	-- 4686: 	lli	%r3, 4
"00010100000000000000000000000000",	-- 4687: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4688: 	lhif	%f0, 0.000000
"00111100010111100000000000000000",	-- 4689: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 4690: 	sw	%r1, [%sp + 1]
"10000100000000110000100000000000",	-- 4691: 	add	%r1, %r0, %r3
"00111111111111100000000000000010",	-- 4692: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 4693: 	addi	%sp, %sp, 3
"01011000000000000010101000100100",	-- 4694: 	jal	yj_create_float_array
"10101011110111100000000000000011",	-- 4695: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 4696: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000000",	-- 4697: 	lli	%r2, 0
"00111011110000110000000000000001",	-- 4698: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4699: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4700: 	lf	%f0, [%r2 + 0]
"00111011110000100000000000000000",	-- 4701: 	lw	%r2, [%sp + 0]
"00111100001111100000000000000010",	-- 4702: 	sw	%r1, [%sp + 2]
"10110000000111100000000000000011",	-- 4703: 	sf	%f0, [%sp + 3]
"10000100000000100000100000000000",	-- 4704: 	add	%r1, %r0, %r2
"00111111111111100000000000000100",	-- 4705: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 4706: 	addi	%sp, %sp, 5
"01011000000000000000011001011010",	-- 4707: 	jal	o_param_a.2632
"10101011110111100000000000000101",	-- 4708: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 4709: 	lw	%ra, [%sp + 4]
"10010011110000010000000000000011",	-- 4710: 	lf	%f1, [%sp + 3]
"11101000001000000000000000000000",	-- 4711: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 4712: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 4713: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 4714: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4715: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4716: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000100",	-- 4717: 	sf	%f0, [%sp + 4]
"10110000001111100000000000000101",	-- 4718: 	sf	%f1, [%sp + 5]
"00111111111111100000000000000110",	-- 4719: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 4720: 	addi	%sp, %sp, 7
"01011000000000000000011001011111",	-- 4721: 	jal	o_param_b.2634
"10101011110111100000000000000111",	-- 4722: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 4723: 	lw	%ra, [%sp + 6]
"10010011110000010000000000000101",	-- 4724: 	lf	%f1, [%sp + 5]
"11101000001000000000000000000000",	-- 4725: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000100",	-- 4726: 	lf	%f1, [%sp + 4]
"11100000001000000000000000000000",	-- 4727: 	addf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 4728: 	lli	%r1, 2
"00111011110000100000000000000001",	-- 4729: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 4730: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4731: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4732: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000110",	-- 4733: 	sf	%f0, [%sp + 6]
"10110000001111100000000000000111",	-- 4734: 	sf	%f1, [%sp + 7]
"00111111111111100000000000001000",	-- 4735: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 4736: 	addi	%sp, %sp, 9
"01011000000000000000011001100100",	-- 4737: 	jal	o_param_c.2636
"10101011110111100000000000001001",	-- 4738: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 4739: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000111",	-- 4740: 	lf	%f1, [%sp + 7]
"11101000001000000000000000000000",	-- 4741: 	mulf	%f0, %f1, %f0
"10010011110000010000000000000110",	-- 4742: 	lf	%f1, [%sp + 6]
"11100000001000000000000000000000",	-- 4743: 	addf	%f0, %f1, %f0
"10110000000111100000000000001000",	-- 4744: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 4745: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4746: 	addi	%sp, %sp, 10
"01011000000000000000010011010110",	-- 4747: 	jal	fispos.2522
"10101011110111100000000000001010",	-- 4748: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4749: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000000",	-- 4750: 	lli	%r2, 0
"00101000001000100000000000001000",	-- 4751: 	bneq	%r1, %r2, bneq_else.9049
"11001100000000010000000000000000",	-- 4752: 	lli	%r1, 0
"00010100000000000000000000000000",	-- 4753: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4754: 	lhif	%f0, 0.000000
"00111011110000100000000000000010",	-- 4755: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4756: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4757: 	sf	%f0, [%r1 + 0]
"01010100000000000001001011011011",	-- 4758: 	j	bneq_cont.9050
	-- bneq_else.9049:
"11001100000000010000000000000000",	-- 4759: 	lli	%r1, 0
"00010100000000000000000000000000",	-- 4760: 	llif	%f0, -1.000000
"00010000000000001011111110000000",	-- 4761: 	lhif	%f0, -1.000000
"10010011110000010000000000001000",	-- 4762: 	lf	%f1, [%sp + 8]
"11101100000000010000000000000000",	-- 4763: 	divf	%f0, %f0, %f1
"00111011110000100000000000000010",	-- 4764: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4765: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4766: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 4767: 	lli	%r1, 1
"00111011110000110000000000000000",	-- 4768: 	lw	%r3, [%sp + 0]
"00111100001111100000000000001001",	-- 4769: 	sw	%r1, [%sp + 9]
"10000100000000110000100000000000",	-- 4770: 	add	%r1, %r0, %r3
"00111111111111100000000000001010",	-- 4771: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4772: 	addi	%sp, %sp, 11
"01011000000000000000011001011010",	-- 4773: 	jal	o_param_a.2632
"10101011110111100000000000001011",	-- 4774: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4775: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001000",	-- 4776: 	lf	%f1, [%sp + 8]
"11101100000000010000000000000000",	-- 4777: 	divf	%f0, %f0, %f1
"00111111111111100000000000001010",	-- 4778: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4779: 	addi	%sp, %sp, 11
"01011000000000000010101001010001",	-- 4780: 	jal	yj_fneg
"10101011110111100000000000001011",	-- 4781: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4782: 	lw	%ra, [%sp + 10]
"00111011110000010000000000001001",	-- 4783: 	lw	%r1, [%sp + 9]
"00111011110000100000000000000010",	-- 4784: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4785: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4786: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 4787: 	lli	%r1, 2
"00111011110000110000000000000000",	-- 4788: 	lw	%r3, [%sp + 0]
"00111100001111100000000000001010",	-- 4789: 	sw	%r1, [%sp + 10]
"10000100000000110000100000000000",	-- 4790: 	add	%r1, %r0, %r3
"00111111111111100000000000001011",	-- 4791: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4792: 	addi	%sp, %sp, 12
"01011000000000000000011001011111",	-- 4793: 	jal	o_param_b.2634
"10101011110111100000000000001100",	-- 4794: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4795: 	lw	%ra, [%sp + 11]
"10010011110000010000000000001000",	-- 4796: 	lf	%f1, [%sp + 8]
"11101100000000010000000000000000",	-- 4797: 	divf	%f0, %f0, %f1
"00111111111111100000000000001011",	-- 4798: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 4799: 	addi	%sp, %sp, 12
"01011000000000000010101001010001",	-- 4800: 	jal	yj_fneg
"10101011110111100000000000001100",	-- 4801: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 4802: 	lw	%ra, [%sp + 11]
"00111011110000010000000000001010",	-- 4803: 	lw	%r1, [%sp + 10]
"00111011110000100000000000000010",	-- 4804: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4805: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4806: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 4807: 	lli	%r1, 3
"00111011110000110000000000000000",	-- 4808: 	lw	%r3, [%sp + 0]
"00111100001111100000000000001011",	-- 4809: 	sw	%r1, [%sp + 11]
"10000100000000110000100000000000",	-- 4810: 	add	%r1, %r0, %r3
"00111111111111100000000000001100",	-- 4811: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4812: 	addi	%sp, %sp, 13
"01011000000000000000011001100100",	-- 4813: 	jal	o_param_c.2636
"10101011110111100000000000001101",	-- 4814: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4815: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001000",	-- 4816: 	lf	%f1, [%sp + 8]
"11101100000000010000000000000000",	-- 4817: 	divf	%f0, %f0, %f1
"00111111111111100000000000001100",	-- 4818: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4819: 	addi	%sp, %sp, 13
"01011000000000000010101001010001",	-- 4820: 	jal	yj_fneg
"10101011110111100000000000001101",	-- 4821: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4822: 	lw	%ra, [%sp + 12]
"00111011110000010000000000001011",	-- 4823: 	lw	%r1, [%sp + 11]
"00111011110000100000000000000010",	-- 4824: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4825: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4826: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9050:
"10000100000000100000100000000000",	-- 4827: 	add	%r1, %r0, %r2
"01001111111000000000000000000000",	-- 4828: 	jr	%ra
	-- setup_second_table.2806:
"11001100000000110000000000000101",	-- 4829: 	lli	%r3, 5
"00010100000000000000000000000000",	-- 4830: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 4831: 	lhif	%f0, 0.000000
"00111100010111100000000000000000",	-- 4832: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 4833: 	sw	%r1, [%sp + 1]
"10000100000000110000100000000000",	-- 4834: 	add	%r1, %r0, %r3
"00111111111111100000000000000010",	-- 4835: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 4836: 	addi	%sp, %sp, 3
"01011000000000000010101000100100",	-- 4837: 	jal	yj_create_float_array
"10101011110111100000000000000011",	-- 4838: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 4839: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000000",	-- 4840: 	lli	%r2, 0
"00111011110000110000000000000001",	-- 4841: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4842: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4843: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000001",	-- 4844: 	lli	%r2, 1
"10000100011000100001000000000000",	-- 4845: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 4846: 	lf	%f1, [%r2 + 0]
"11001100000000100000000000000010",	-- 4847: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 4848: 	add	%r2, %r3, %r2
"10010000010000100000000000000000",	-- 4849: 	lf	%f2, [%r2 + 0]
"00111011110000100000000000000000",	-- 4850: 	lw	%r2, [%sp + 0]
"00111100001111100000000000000010",	-- 4851: 	sw	%r1, [%sp + 2]
"10000100000000100000100000000000",	-- 4852: 	add	%r1, %r0, %r2
"00111111111111100000000000000011",	-- 4853: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 4854: 	addi	%sp, %sp, 4
"01011000000000000000110001111010",	-- 4855: 	jal	quadratic.2737
"10101011110111100000000000000100",	-- 4856: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 4857: 	lw	%ra, [%sp + 3]
"11001100000000010000000000000000",	-- 4858: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 4859: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 4860: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4861: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4862: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000011",	-- 4863: 	sf	%f0, [%sp + 3]
"10110000001111100000000000000100",	-- 4864: 	sf	%f1, [%sp + 4]
"00111111111111100000000000000101",	-- 4865: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 4866: 	addi	%sp, %sp, 6
"01011000000000000000011001011010",	-- 4867: 	jal	o_param_a.2632
"10101011110111100000000000000110",	-- 4868: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 4869: 	lw	%ra, [%sp + 5]
"10010011110000010000000000000100",	-- 4870: 	lf	%f1, [%sp + 4]
"11101000001000000000000000000000",	-- 4871: 	mulf	%f0, %f1, %f0
"00111111111111100000000000000101",	-- 4872: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 4873: 	addi	%sp, %sp, 6
"01011000000000000010101001010001",	-- 4874: 	jal	yj_fneg
"10101011110111100000000000000110",	-- 4875: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 4876: 	lw	%ra, [%sp + 5]
"11001100000000010000000000000001",	-- 4877: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 4878: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 4879: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4880: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4881: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000101",	-- 4882: 	sf	%f0, [%sp + 5]
"10110000001111100000000000000110",	-- 4883: 	sf	%f1, [%sp + 6]
"00111111111111100000000000000111",	-- 4884: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 4885: 	addi	%sp, %sp, 8
"01011000000000000000011001011111",	-- 4886: 	jal	o_param_b.2634
"10101011110111100000000000001000",	-- 4887: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 4888: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000110",	-- 4889: 	lf	%f1, [%sp + 6]
"11101000001000000000000000000000",	-- 4890: 	mulf	%f0, %f1, %f0
"00111111111111100000000000000111",	-- 4891: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 4892: 	addi	%sp, %sp, 8
"01011000000000000010101001010001",	-- 4893: 	jal	yj_fneg
"10101011110111100000000000001000",	-- 4894: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 4895: 	lw	%ra, [%sp + 7]
"11001100000000010000000000000010",	-- 4896: 	lli	%r1, 2
"00111011110000100000000000000001",	-- 4897: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 4898: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4899: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4900: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000111",	-- 4901: 	sf	%f0, [%sp + 7]
"10110000001111100000000000001000",	-- 4902: 	sf	%f1, [%sp + 8]
"00111111111111100000000000001001",	-- 4903: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4904: 	addi	%sp, %sp, 10
"01011000000000000000011001100100",	-- 4905: 	jal	o_param_c.2636
"10101011110111100000000000001010",	-- 4906: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4907: 	lw	%ra, [%sp + 9]
"10010011110000010000000000001000",	-- 4908: 	lf	%f1, [%sp + 8]
"11101000001000000000000000000000",	-- 4909: 	mulf	%f0, %f1, %f0
"00111111111111100000000000001001",	-- 4910: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 4911: 	addi	%sp, %sp, 10
"01011000000000000010101001010001",	-- 4912: 	jal	yj_fneg
"10101011110111100000000000001010",	-- 4913: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 4914: 	lw	%ra, [%sp + 9]
"11001100000000010000000000000000",	-- 4915: 	lli	%r1, 0
"00111011110000100000000000000010",	-- 4916: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4917: 	add	%r1, %r2, %r1
"10010011110000010000000000000011",	-- 4918: 	lf	%f1, [%sp + 3]
"10110000001000010000000000000000",	-- 4919: 	sf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4920: 	lw	%r1, [%sp + 0]
"10110000000111100000000000001001",	-- 4921: 	sf	%f0, [%sp + 9]
"00111111111111100000000000001010",	-- 4922: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 4923: 	addi	%sp, %sp, 11
"01011000000000000000011001011000",	-- 4924: 	jal	o_isrot.2630
"10101011110111100000000000001011",	-- 4925: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 4926: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 4927: 	lli	%r2, 0
"00101000001000100000000000001111",	-- 4928: 	bneq	%r1, %r2, bneq_else.9051
"11001100000000010000000000000001",	-- 4929: 	lli	%r1, 1
"00111011110000100000000000000010",	-- 4930: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4931: 	add	%r1, %r2, %r1
"10010011110000000000000000000101",	-- 4932: 	lf	%f0, [%sp + 5]
"10110000000000010000000000000000",	-- 4933: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 4934: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 4935: 	add	%r1, %r2, %r1
"10010011110000000000000000000111",	-- 4936: 	lf	%f0, [%sp + 7]
"10110000000000010000000000000000",	-- 4937: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 4938: 	lli	%r1, 3
"10000100010000010000100000000000",	-- 4939: 	add	%r1, %r2, %r1
"10010011110000000000000000001001",	-- 4940: 	lf	%f0, [%sp + 9]
"10110000000000010000000000000000",	-- 4941: 	sf	%f0, [%r1 + 0]
"01010100000000000001001111010000",	-- 4942: 	j	bneq_cont.9052
	-- bneq_else.9051:
"11001100000000010000000000000001",	-- 4943: 	lli	%r1, 1
"11001100000000100000000000000010",	-- 4944: 	lli	%r2, 2
"00111011110000110000000000000001",	-- 4945: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 4946: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 4947: 	lf	%f0, [%r2 + 0]
"00111011110000100000000000000000",	-- 4948: 	lw	%r2, [%sp + 0]
"00111100001111100000000000001010",	-- 4949: 	sw	%r1, [%sp + 10]
"10110000000111100000000000001011",	-- 4950: 	sf	%f0, [%sp + 11]
"10000100000000100000100000000000",	-- 4951: 	add	%r1, %r0, %r2
"00111111111111100000000000001100",	-- 4952: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 4953: 	addi	%sp, %sp, 13
"01011000000000000000011010011000",	-- 4954: 	jal	o_param_r2.2658
"10101011110111100000000000001101",	-- 4955: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 4956: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001011",	-- 4957: 	lf	%f1, [%sp + 11]
"11101000001000000000000000000000",	-- 4958: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 4959: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 4960: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 4961: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 4962: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 4963: 	lw	%r1, [%sp + 0]
"10110000000111100000000000001100",	-- 4964: 	sf	%f0, [%sp + 12]
"10110000001111100000000000001101",	-- 4965: 	sf	%f1, [%sp + 13]
"00111111111111100000000000001110",	-- 4966: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 4967: 	addi	%sp, %sp, 15
"01011000000000000000011010011101",	-- 4968: 	jal	o_param_r3.2660
"10101011110111100000000000001111",	-- 4969: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 4970: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001101",	-- 4971: 	lf	%f1, [%sp + 13]
"11101000001000000000000000000000",	-- 4972: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001100",	-- 4973: 	lf	%f1, [%sp + 12]
"11100000001000000000000000000000",	-- 4974: 	addf	%f0, %f1, %f0
"00111111111111100000000000001110",	-- 4975: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 4976: 	addi	%sp, %sp, 15
"01011000000000000000010011101101",	-- 4977: 	jal	fhalf.2528
"10101011110111100000000000001111",	-- 4978: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 4979: 	lw	%ra, [%sp + 14]
"10010011110000010000000000000101",	-- 4980: 	lf	%f1, [%sp + 5]
"11100100001000000000000000000000",	-- 4981: 	subf	%f0, %f1, %f0
"00111011110000010000000000001010",	-- 4982: 	lw	%r1, [%sp + 10]
"00111011110000100000000000000010",	-- 4983: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 4984: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 4985: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 4986: 	lli	%r1, 2
"11001100000000110000000000000010",	-- 4987: 	lli	%r3, 2
"00111011110001000000000000000001",	-- 4988: 	lw	%r4, [%sp + 1]
"10000100100000110001100000000000",	-- 4989: 	add	%r3, %r4, %r3
"10010000011000000000000000000000",	-- 4990: 	lf	%f0, [%r3 + 0]
"00111011110000110000000000000000",	-- 4991: 	lw	%r3, [%sp + 0]
"00111100001111100000000000001110",	-- 4992: 	sw	%r1, [%sp + 14]
"10110000000111100000000000001111",	-- 4993: 	sf	%f0, [%sp + 15]
"10000100000000110000100000000000",	-- 4994: 	add	%r1, %r0, %r3
"00111111111111100000000000010000",	-- 4995: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 4996: 	addi	%sp, %sp, 17
"01011000000000000000011010010011",	-- 4997: 	jal	o_param_r1.2656
"10101011110111100000000000010001",	-- 4998: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 4999: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001111",	-- 5000: 	lf	%f1, [%sp + 15]
"11101000001000000000000000000000",	-- 5001: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 5002: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 5003: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 5004: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 5005: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 5006: 	lw	%r1, [%sp + 0]
"10110000000111100000000000010000",	-- 5007: 	sf	%f0, [%sp + 16]
"10110000001111100000000000010001",	-- 5008: 	sf	%f1, [%sp + 17]
"00111111111111100000000000010010",	-- 5009: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 5010: 	addi	%sp, %sp, 19
"01011000000000000000011010011101",	-- 5011: 	jal	o_param_r3.2660
"10101011110111100000000000010011",	-- 5012: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 5013: 	lw	%ra, [%sp + 18]
"10010011110000010000000000010001",	-- 5014: 	lf	%f1, [%sp + 17]
"11101000001000000000000000000000",	-- 5015: 	mulf	%f0, %f1, %f0
"10010011110000010000000000010000",	-- 5016: 	lf	%f1, [%sp + 16]
"11100000001000000000000000000000",	-- 5017: 	addf	%f0, %f1, %f0
"00111111111111100000000000010010",	-- 5018: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 5019: 	addi	%sp, %sp, 19
"01011000000000000000010011101101",	-- 5020: 	jal	fhalf.2528
"10101011110111100000000000010011",	-- 5021: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 5022: 	lw	%ra, [%sp + 18]
"10010011110000010000000000000111",	-- 5023: 	lf	%f1, [%sp + 7]
"11100100001000000000000000000000",	-- 5024: 	subf	%f0, %f1, %f0
"00111011110000010000000000001110",	-- 5025: 	lw	%r1, [%sp + 14]
"00111011110000100000000000000010",	-- 5026: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 5027: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5028: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000011",	-- 5029: 	lli	%r1, 3
"11001100000000110000000000000001",	-- 5030: 	lli	%r3, 1
"00111011110001000000000000000001",	-- 5031: 	lw	%r4, [%sp + 1]
"10000100100000110001100000000000",	-- 5032: 	add	%r3, %r4, %r3
"10010000011000000000000000000000",	-- 5033: 	lf	%f0, [%r3 + 0]
"00111011110000110000000000000000",	-- 5034: 	lw	%r3, [%sp + 0]
"00111100001111100000000000010010",	-- 5035: 	sw	%r1, [%sp + 18]
"10110000000111100000000000010011",	-- 5036: 	sf	%f0, [%sp + 19]
"10000100000000110000100000000000",	-- 5037: 	add	%r1, %r0, %r3
"00111111111111100000000000010100",	-- 5038: 	sw	%ra, [%sp + 20]
"10100111110111100000000000010101",	-- 5039: 	addi	%sp, %sp, 21
"01011000000000000000011010010011",	-- 5040: 	jal	o_param_r1.2656
"10101011110111100000000000010101",	-- 5041: 	subi	%sp, %sp, 21
"00111011110111110000000000010100",	-- 5042: 	lw	%ra, [%sp + 20]
"10010011110000010000000000010011",	-- 5043: 	lf	%f1, [%sp + 19]
"11101000001000000000000000000000",	-- 5044: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 5045: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 5046: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 5047: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 5048: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000000",	-- 5049: 	lw	%r1, [%sp + 0]
"10110000000111100000000000010100",	-- 5050: 	sf	%f0, [%sp + 20]
"10110000001111100000000000010101",	-- 5051: 	sf	%f1, [%sp + 21]
"00111111111111100000000000010110",	-- 5052: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 5053: 	addi	%sp, %sp, 23
"01011000000000000000011010011000",	-- 5054: 	jal	o_param_r2.2658
"10101011110111100000000000010111",	-- 5055: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 5056: 	lw	%ra, [%sp + 22]
"10010011110000010000000000010101",	-- 5057: 	lf	%f1, [%sp + 21]
"11101000001000000000000000000000",	-- 5058: 	mulf	%f0, %f1, %f0
"10010011110000010000000000010100",	-- 5059: 	lf	%f1, [%sp + 20]
"11100000001000000000000000000000",	-- 5060: 	addf	%f0, %f1, %f0
"00111111111111100000000000010110",	-- 5061: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 5062: 	addi	%sp, %sp, 23
"01011000000000000000010011101101",	-- 5063: 	jal	fhalf.2528
"10101011110111100000000000010111",	-- 5064: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 5065: 	lw	%ra, [%sp + 22]
"10010011110000010000000000001001",	-- 5066: 	lf	%f1, [%sp + 9]
"11100100001000000000000000000000",	-- 5067: 	subf	%f0, %f1, %f0
"00111011110000010000000000010010",	-- 5068: 	lw	%r1, [%sp + 18]
"00111011110000100000000000000010",	-- 5069: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 5070: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5071: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9052:
"10010011110000000000000000000011",	-- 5072: 	lf	%f0, [%sp + 3]
"00111111111111100000000000010110",	-- 5073: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 5074: 	addi	%sp, %sp, 23
"01011000000000000000010011100100",	-- 5075: 	jal	fiszero.2526
"10101011110111100000000000010111",	-- 5076: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 5077: 	lw	%ra, [%sp + 22]
"11001100000000100000000000000000",	-- 5078: 	lli	%r2, 0
"00101000001000100000000000001010",	-- 5079: 	bneq	%r1, %r2, bneq_else.9053
"11001100000000010000000000000100",	-- 5080: 	lli	%r1, 4
"00010100000000000000000000000000",	-- 5081: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 5082: 	lhif	%f0, 1.000000
"10010011110000010000000000000011",	-- 5083: 	lf	%f1, [%sp + 3]
"11101100000000010000000000000000",	-- 5084: 	divf	%f0, %f0, %f1
"00111011110000100000000000000010",	-- 5085: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 5086: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5087: 	sf	%f0, [%r1 + 0]
"01010100000000000001001111100001",	-- 5088: 	j	bneq_cont.9054
	-- bneq_else.9053:
	-- bneq_cont.9054:
"00111011110000010000000000000010",	-- 5089: 	lw	%r1, [%sp + 2]
"01001111111000000000000000000000",	-- 5090: 	jr	%ra
	-- iter_setup_dirvec_constants.2809:
"00111011011000110000000000000001",	-- 5091: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 5092: 	lli	%r4, 0
"00110000100000100000000001001001",	-- 5093: 	bgt	%r4, %r2, bgt_else.9055
"10000100011000100001100000000000",	-- 5094: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 5095: 	lw	%r3, [%r3 + 0]
"00111111011111100000000000000000",	-- 5096: 	sw	%r27, [%sp + 0]
"00111100010111100000000000000001",	-- 5097: 	sw	%r2, [%sp + 1]
"00111100011111100000000000000010",	-- 5098: 	sw	%r3, [%sp + 2]
"00111100001111100000000000000011",	-- 5099: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 5100: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5101: 	addi	%sp, %sp, 5
"01011000000000000000011010111110",	-- 5102: 	jal	d_const.2685
"10101011110111100000000000000101",	-- 5103: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5104: 	lw	%ra, [%sp + 4]
"00111011110000100000000000000011",	-- 5105: 	lw	%r2, [%sp + 3]
"00111100001111100000000000000100",	-- 5106: 	sw	%r1, [%sp + 4]
"10000100000000100000100000000000",	-- 5107: 	add	%r1, %r0, %r2
"00111111111111100000000000000101",	-- 5108: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5109: 	addi	%sp, %sp, 6
"01011000000000000000011010111100",	-- 5110: 	jal	d_vec.2683
"10101011110111100000000000000110",	-- 5111: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5112: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000010",	-- 5113: 	lw	%r2, [%sp + 2]
"00111100001111100000000000000101",	-- 5114: 	sw	%r1, [%sp + 5]
"10000100000000100000100000000000",	-- 5115: 	add	%r1, %r0, %r2
"00111111111111100000000000000110",	-- 5116: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5117: 	addi	%sp, %sp, 7
"01011000000000000000011001010010",	-- 5118: 	jal	o_form.2624
"10101011110111100000000000000111",	-- 5119: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5120: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000001",	-- 5121: 	lli	%r2, 1
"00101000001000100000000000001101",	-- 5122: 	bneq	%r1, %r2, bneq_else.9056
"00111011110000010000000000000101",	-- 5123: 	lw	%r1, [%sp + 5]
"00111011110000100000000000000010",	-- 5124: 	lw	%r2, [%sp + 2]
"00111111111111100000000000000110",	-- 5125: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5126: 	addi	%sp, %sp, 7
"01011000000000000001000101101000",	-- 5127: 	jal	setup_rect_table.2800
"10101011110111100000000000000111",	-- 5128: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5129: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000001",	-- 5130: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000100",	-- 5131: 	lw	%r3, [%sp + 4]
"10000100011000100001100000000000",	-- 5132: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 5133: 	sw	%r1, [%r3 + 0]
"01010100000000000001010000101000",	-- 5134: 	j	bneq_cont.9057
	-- bneq_else.9056:
"11001100000000100000000000000010",	-- 5135: 	lli	%r2, 2
"00101000001000100000000000001101",	-- 5136: 	bneq	%r1, %r2, bneq_else.9058
"00111011110000010000000000000101",	-- 5137: 	lw	%r1, [%sp + 5]
"00111011110000100000000000000010",	-- 5138: 	lw	%r2, [%sp + 2]
"00111111111111100000000000000110",	-- 5139: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5140: 	addi	%sp, %sp, 7
"01011000000000000001001001001110",	-- 5141: 	jal	setup_surface_table.2803
"10101011110111100000000000000111",	-- 5142: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5143: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000001",	-- 5144: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000100",	-- 5145: 	lw	%r3, [%sp + 4]
"10000100011000100001100000000000",	-- 5146: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 5147: 	sw	%r1, [%r3 + 0]
"01010100000000000001010000101000",	-- 5148: 	j	bneq_cont.9059
	-- bneq_else.9058:
"00111011110000010000000000000101",	-- 5149: 	lw	%r1, [%sp + 5]
"00111011110000100000000000000010",	-- 5150: 	lw	%r2, [%sp + 2]
"00111111111111100000000000000110",	-- 5151: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5152: 	addi	%sp, %sp, 7
"01011000000000000001001011011101",	-- 5153: 	jal	setup_second_table.2806
"10101011110111100000000000000111",	-- 5154: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5155: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000001",	-- 5156: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000100",	-- 5157: 	lw	%r3, [%sp + 4]
"10000100011000100001100000000000",	-- 5158: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 5159: 	sw	%r1, [%r3 + 0]
	-- bneq_cont.9059:
	-- bneq_cont.9057:
"11001100000000010000000000000001",	-- 5160: 	lli	%r1, 1
"10001000010000010001000000000000",	-- 5161: 	sub	%r2, %r2, %r1
"00111011110000010000000000000011",	-- 5162: 	lw	%r1, [%sp + 3]
"00111011110110110000000000000000",	-- 5163: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 5164: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5165: 	jr	%r26
	-- bgt_else.9055:
"01001111111000000000000000000000",	-- 5166: 	jr	%ra
	-- setup_dirvec_constants.2812:
"00111011011000100000000000000010",	-- 5167: 	lw	%r2, [%r27 + 2]
"00111011011110110000000000000001",	-- 5168: 	lw	%r27, [%r27 + 1]
"11001100000000110000000000000000",	-- 5169: 	lli	%r3, 0
"10000100010000110001000000000000",	-- 5170: 	add	%r2, %r2, %r3
"00111000010000100000000000000000",	-- 5171: 	lw	%r2, [%r2 + 0]
"11001100000000110000000000000001",	-- 5172: 	lli	%r3, 1
"10001000010000110001000000000000",	-- 5173: 	sub	%r2, %r2, %r3
"00111011011110100000000000000000",	-- 5174: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5175: 	jr	%r26
	-- setup_startp_constants.2814:
"00111011011000110000000000000001",	-- 5176: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 5177: 	lli	%r4, 0
"00110000100000100000000010010110",	-- 5178: 	bgt	%r4, %r2, bgt_else.9061
"10000100011000100001100000000000",	-- 5179: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 5180: 	lw	%r3, [%r3 + 0]
"00111111011111100000000000000000",	-- 5181: 	sw	%r27, [%sp + 0]
"00111100010111100000000000000001",	-- 5182: 	sw	%r2, [%sp + 1]
"00111100001111100000000000000010",	-- 5183: 	sw	%r1, [%sp + 2]
"00111100011111100000000000000011",	-- 5184: 	sw	%r3, [%sp + 3]
"10000100000000110000100000000000",	-- 5185: 	add	%r1, %r0, %r3
"00111111111111100000000000000100",	-- 5186: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5187: 	addi	%sp, %sp, 5
"01011000000000000000011010100010",	-- 5188: 	jal	o_param_ctbl.2662
"10101011110111100000000000000101",	-- 5189: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5190: 	lw	%ra, [%sp + 4]
"00111011110000100000000000000011",	-- 5191: 	lw	%r2, [%sp + 3]
"00111100001111100000000000000100",	-- 5192: 	sw	%r1, [%sp + 4]
"10000100000000100000100000000000",	-- 5193: 	add	%r1, %r0, %r2
"00111111111111100000000000000101",	-- 5194: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5195: 	addi	%sp, %sp, 6
"01011000000000000000011001010010",	-- 5196: 	jal	o_form.2624
"10101011110111100000000000000110",	-- 5197: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5198: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000000",	-- 5199: 	lli	%r2, 0
"11001100000000110000000000000000",	-- 5200: 	lli	%r3, 0
"00111011110001000000000000000010",	-- 5201: 	lw	%r4, [%sp + 2]
"10000100100000110001100000000000",	-- 5202: 	add	%r3, %r4, %r3
"10010000011000000000000000000000",	-- 5203: 	lf	%f0, [%r3 + 0]
"00111011110000110000000000000011",	-- 5204: 	lw	%r3, [%sp + 3]
"00111100001111100000000000000101",	-- 5205: 	sw	%r1, [%sp + 5]
"00111100010111100000000000000110",	-- 5206: 	sw	%r2, [%sp + 6]
"10110000000111100000000000000111",	-- 5207: 	sf	%f0, [%sp + 7]
"10000100000000110000100000000000",	-- 5208: 	add	%r1, %r0, %r3
"00111111111111100000000000001000",	-- 5209: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 5210: 	addi	%sp, %sp, 9
"01011000000000000000011001101011",	-- 5211: 	jal	o_param_x.2640
"10101011110111100000000000001001",	-- 5212: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 5213: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000111",	-- 5214: 	lf	%f1, [%sp + 7]
"11100100001000000000000000000000",	-- 5215: 	subf	%f0, %f1, %f0
"00111011110000010000000000000110",	-- 5216: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000100",	-- 5217: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5218: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5219: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 5220: 	lli	%r1, 1
"11001100000000110000000000000001",	-- 5221: 	lli	%r3, 1
"00111011110001000000000000000010",	-- 5222: 	lw	%r4, [%sp + 2]
"10000100100000110001100000000000",	-- 5223: 	add	%r3, %r4, %r3
"10010000011000000000000000000000",	-- 5224: 	lf	%f0, [%r3 + 0]
"00111011110000110000000000000011",	-- 5225: 	lw	%r3, [%sp + 3]
"00111100001111100000000000001000",	-- 5226: 	sw	%r1, [%sp + 8]
"10110000000111100000000000001001",	-- 5227: 	sf	%f0, [%sp + 9]
"10000100000000110000100000000000",	-- 5228: 	add	%r1, %r0, %r3
"00111111111111100000000000001010",	-- 5229: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 5230: 	addi	%sp, %sp, 11
"01011000000000000000011001110000",	-- 5231: 	jal	o_param_y.2642
"10101011110111100000000000001011",	-- 5232: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 5233: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 5234: 	lf	%f1, [%sp + 9]
"11100100001000000000000000000000",	-- 5235: 	subf	%f0, %f1, %f0
"00111011110000010000000000001000",	-- 5236: 	lw	%r1, [%sp + 8]
"00111011110000100000000000000100",	-- 5237: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5238: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5239: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 5240: 	lli	%r1, 2
"11001100000000110000000000000010",	-- 5241: 	lli	%r3, 2
"00111011110001000000000000000010",	-- 5242: 	lw	%r4, [%sp + 2]
"10000100100000110001100000000000",	-- 5243: 	add	%r3, %r4, %r3
"10010000011000000000000000000000",	-- 5244: 	lf	%f0, [%r3 + 0]
"00111011110000110000000000000011",	-- 5245: 	lw	%r3, [%sp + 3]
"00111100001111100000000000001010",	-- 5246: 	sw	%r1, [%sp + 10]
"10110000000111100000000000001011",	-- 5247: 	sf	%f0, [%sp + 11]
"10000100000000110000100000000000",	-- 5248: 	add	%r1, %r0, %r3
"00111111111111100000000000001100",	-- 5249: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 5250: 	addi	%sp, %sp, 13
"01011000000000000000011001110101",	-- 5251: 	jal	o_param_z.2644
"10101011110111100000000000001101",	-- 5252: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 5253: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001011",	-- 5254: 	lf	%f1, [%sp + 11]
"11100100001000000000000000000000",	-- 5255: 	subf	%f0, %f1, %f0
"00111011110000010000000000001010",	-- 5256: 	lw	%r1, [%sp + 10]
"00111011110000100000000000000100",	-- 5257: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5258: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5259: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 5260: 	lli	%r1, 2
"00111011110000110000000000000101",	-- 5261: 	lw	%r3, [%sp + 5]
"00101000011000010000000000011110",	-- 5262: 	bneq	%r3, %r1, bneq_else.9062
"11001100000000010000000000000011",	-- 5263: 	lli	%r1, 3
"00111011110000110000000000000011",	-- 5264: 	lw	%r3, [%sp + 3]
"00111100001111100000000000001100",	-- 5265: 	sw	%r1, [%sp + 12]
"10000100000000110000100000000000",	-- 5266: 	add	%r1, %r0, %r3
"00111111111111100000000000001101",	-- 5267: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 5268: 	addi	%sp, %sp, 14
"01011000000000000000011001101001",	-- 5269: 	jal	o_param_abc.2638
"10101011110111100000000000001110",	-- 5270: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 5271: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 5272: 	lli	%r2, 0
"00111011110000110000000000000100",	-- 5273: 	lw	%r3, [%sp + 4]
"10000100011000100001000000000000",	-- 5274: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 5275: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000001",	-- 5276: 	lli	%r2, 1
"10000100011000100001000000000000",	-- 5277: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 5278: 	lf	%f1, [%r2 + 0]
"11001100000000100000000000000010",	-- 5279: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 5280: 	add	%r2, %r3, %r2
"10010000010000100000000000000000",	-- 5281: 	lf	%f2, [%r2 + 0]
"00111111111111100000000000001101",	-- 5282: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 5283: 	addi	%sp, %sp, 14
"01011000000000000000010110111111",	-- 5284: 	jal	veciprod2.2600
"10101011110111100000000000001110",	-- 5285: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 5286: 	lw	%ra, [%sp + 13]
"00111011110000010000000000001100",	-- 5287: 	lw	%r1, [%sp + 12]
"00111011110000100000000000000100",	-- 5288: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5289: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5290: 	sf	%f0, [%r1 + 0]
"01010100000000000001010011001001",	-- 5291: 	j	bneq_cont.9063
	-- bneq_else.9062:
"11001100000000010000000000000010",	-- 5292: 	lli	%r1, 2
"00110000011000010000000000000010",	-- 5293: 	bgt	%r3, %r1, bgt_else.9064
"01010100000000000001010011001001",	-- 5294: 	j	bgt_cont.9065
	-- bgt_else.9064:
"11001100000000010000000000000000",	-- 5295: 	lli	%r1, 0
"10000100010000010000100000000000",	-- 5296: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 5297: 	lf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 5298: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 5299: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 5300: 	lf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 5301: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 5302: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 5303: 	lf	%f2, [%r1 + 0]
"00111011110000010000000000000011",	-- 5304: 	lw	%r1, [%sp + 3]
"00111111111111100000000000001101",	-- 5305: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 5306: 	addi	%sp, %sp, 14
"01011000000000000000110001111010",	-- 5307: 	jal	quadratic.2737
"10101011110111100000000000001110",	-- 5308: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 5309: 	lw	%ra, [%sp + 13]
"11001100000000010000000000000011",	-- 5310: 	lli	%r1, 3
"11001100000000100000000000000011",	-- 5311: 	lli	%r2, 3
"00111011110000110000000000000101",	-- 5312: 	lw	%r3, [%sp + 5]
"00101000011000100000000000000101",	-- 5313: 	bneq	%r3, %r2, bneq_else.9066
"00010100000000010000000000000000",	-- 5314: 	llif	%f1, 1.000000
"00010000000000010011111110000000",	-- 5315: 	lhif	%f1, 1.000000
"11100100000000010000000000000000",	-- 5316: 	subf	%f0, %f0, %f1
"01010100000000000001010011000110",	-- 5317: 	j	bneq_cont.9067
	-- bneq_else.9066:
	-- bneq_cont.9067:
"00111011110000100000000000000100",	-- 5318: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5319: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 5320: 	sf	%f0, [%r1 + 0]
	-- bgt_cont.9065:
	-- bneq_cont.9063:
"11001100000000010000000000000001",	-- 5321: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 5322: 	lw	%r2, [%sp + 1]
"10001000010000010001000000000000",	-- 5323: 	sub	%r2, %r2, %r1
"00111011110000010000000000000010",	-- 5324: 	lw	%r1, [%sp + 2]
"00111011110110110000000000000000",	-- 5325: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 5326: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5327: 	jr	%r26
	-- bgt_else.9061:
"01001111111000000000000000000000",	-- 5328: 	jr	%ra
	-- setup_startp.2817:
"00111011011000100000000000000011",	-- 5329: 	lw	%r2, [%r27 + 3]
"00111011011000110000000000000010",	-- 5330: 	lw	%r3, [%r27 + 2]
"00111011011001000000000000000001",	-- 5331: 	lw	%r4, [%r27 + 1]
"00111100001111100000000000000000",	-- 5332: 	sw	%r1, [%sp + 0]
"00111100011111100000000000000001",	-- 5333: 	sw	%r3, [%sp + 1]
"00111100100111100000000000000010",	-- 5334: 	sw	%r4, [%sp + 2]
"10000100000000101101000000000000",	-- 5335: 	add	%r26, %r0, %r2
"10000100000000010001000000000000",	-- 5336: 	add	%r2, %r0, %r1
"10000100000110100000100000000000",	-- 5337: 	add	%r1, %r0, %r26
"00111111111111100000000000000011",	-- 5338: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 5339: 	addi	%sp, %sp, 4
"01011000000000000000010100111101",	-- 5340: 	jal	veccpy.2586
"10101011110111100000000000000100",	-- 5341: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 5342: 	lw	%ra, [%sp + 3]
"11001100000000010000000000000000",	-- 5343: 	lli	%r1, 0
"00111011110000100000000000000010",	-- 5344: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 5345: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 5346: 	lw	%r1, [%r1 + 0]
"11001100000000100000000000000001",	-- 5347: 	lli	%r2, 1
"10001000001000100001000000000000",	-- 5348: 	sub	%r2, %r1, %r2
"00111011110000010000000000000000",	-- 5349: 	lw	%r1, [%sp + 0]
"00111011110110110000000000000001",	-- 5350: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 5351: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5352: 	jr	%r26
	-- is_rect_outside.2819:
"10110000010111100000000000000000",	-- 5353: 	sf	%f2, [%sp + 0]
"10110000001111100000000000000001",	-- 5354: 	sf	%f1, [%sp + 1]
"00111100001111100000000000000010",	-- 5355: 	sw	%r1, [%sp + 2]
"00111111111111100000000000000011",	-- 5356: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 5357: 	addi	%sp, %sp, 4
"01011000000000000010101001001111",	-- 5358: 	jal	yj_fabs
"10101011110111100000000000000100",	-- 5359: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 5360: 	lw	%ra, [%sp + 3]
"00111011110000010000000000000010",	-- 5361: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000011",	-- 5362: 	sf	%f0, [%sp + 3]
"00111111111111100000000000000100",	-- 5363: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5364: 	addi	%sp, %sp, 5
"01011000000000000000011001011010",	-- 5365: 	jal	o_param_a.2632
"10101011110111100000000000000101",	-- 5366: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5367: 	lw	%ra, [%sp + 4]
"00001100000000010000000000000000",	-- 5368: 	movf	%f1, %f0
"10010011110000000000000000000011",	-- 5369: 	lf	%f0, [%sp + 3]
"00111111111111100000000000000100",	-- 5370: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5371: 	addi	%sp, %sp, 5
"01011000000000000000010011110011",	-- 5372: 	jal	fless.2532
"10101011110111100000000000000101",	-- 5373: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5374: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000000",	-- 5375: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5376: 	bneq	%r1, %r2, bneq_else.9069
"11001100000000010000000000000000",	-- 5377: 	lli	%r1, 0
"01010100000000000001010100101111",	-- 5378: 	j	bneq_cont.9070
	-- bneq_else.9069:
"10010011110000000000000000000001",	-- 5379: 	lf	%f0, [%sp + 1]
"00111111111111100000000000000100",	-- 5380: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5381: 	addi	%sp, %sp, 5
"01011000000000000010101001001111",	-- 5382: 	jal	yj_fabs
"10101011110111100000000000000101",	-- 5383: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5384: 	lw	%ra, [%sp + 4]
"00111011110000010000000000000010",	-- 5385: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000100",	-- 5386: 	sf	%f0, [%sp + 4]
"00111111111111100000000000000101",	-- 5387: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5388: 	addi	%sp, %sp, 6
"01011000000000000000011001011111",	-- 5389: 	jal	o_param_b.2634
"10101011110111100000000000000110",	-- 5390: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5391: 	lw	%ra, [%sp + 5]
"00001100000000010000000000000000",	-- 5392: 	movf	%f1, %f0
"10010011110000000000000000000100",	-- 5393: 	lf	%f0, [%sp + 4]
"00111111111111100000000000000101",	-- 5394: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5395: 	addi	%sp, %sp, 6
"01011000000000000000010011110011",	-- 5396: 	jal	fless.2532
"10101011110111100000000000000110",	-- 5397: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5398: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000000",	-- 5399: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5400: 	bneq	%r1, %r2, bneq_else.9071
"11001100000000010000000000000000",	-- 5401: 	lli	%r1, 0
"01010100000000000001010100101111",	-- 5402: 	j	bneq_cont.9072
	-- bneq_else.9071:
"10010011110000000000000000000000",	-- 5403: 	lf	%f0, [%sp + 0]
"00111111111111100000000000000101",	-- 5404: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5405: 	addi	%sp, %sp, 6
"01011000000000000010101001001111",	-- 5406: 	jal	yj_fabs
"10101011110111100000000000000110",	-- 5407: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5408: 	lw	%ra, [%sp + 5]
"00111011110000010000000000000010",	-- 5409: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000101",	-- 5410: 	sf	%f0, [%sp + 5]
"00111111111111100000000000000110",	-- 5411: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5412: 	addi	%sp, %sp, 7
"01011000000000000000011001100100",	-- 5413: 	jal	o_param_c.2636
"10101011110111100000000000000111",	-- 5414: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5415: 	lw	%ra, [%sp + 6]
"00001100000000010000000000000000",	-- 5416: 	movf	%f1, %f0
"10010011110000000000000000000101",	-- 5417: 	lf	%f0, [%sp + 5]
"00111111111111100000000000000110",	-- 5418: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5419: 	addi	%sp, %sp, 7
"01011000000000000000010011110011",	-- 5420: 	jal	fless.2532
"10101011110111100000000000000111",	-- 5421: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5422: 	lw	%ra, [%sp + 6]
	-- bneq_cont.9072:
	-- bneq_cont.9070:
"11001100000000100000000000000000",	-- 5423: 	lli	%r2, 0
"00101000001000100000000000001101",	-- 5424: 	bneq	%r1, %r2, bneq_else.9073
"00111011110000010000000000000010",	-- 5425: 	lw	%r1, [%sp + 2]
"00111111111111100000000000000110",	-- 5426: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5427: 	addi	%sp, %sp, 7
"01011000000000000000011001010110",	-- 5428: 	jal	o_isinvert.2628
"10101011110111100000000000000111",	-- 5429: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5430: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5431: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5432: 	bneq	%r1, %r2, bneq_else.9074
"11001100000000010000000000000001",	-- 5433: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5434: 	jr	%ra
	-- bneq_else.9074:
"11001100000000010000000000000000",	-- 5435: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5436: 	jr	%ra
	-- bneq_else.9073:
"00111011110000010000000000000010",	-- 5437: 	lw	%r1, [%sp + 2]
"01010100000000000000011001010110",	-- 5438: 	j	o_isinvert.2628
	-- is_plane_outside.2824:
"00111100001111100000000000000000",	-- 5439: 	sw	%r1, [%sp + 0]
"10110000010111100000000000000001",	-- 5440: 	sf	%f2, [%sp + 1]
"10110000001111100000000000000010",	-- 5441: 	sf	%f1, [%sp + 2]
"10110000000111100000000000000011",	-- 5442: 	sf	%f0, [%sp + 3]
"00111111111111100000000000000100",	-- 5443: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5444: 	addi	%sp, %sp, 5
"01011000000000000000011001101001",	-- 5445: 	jal	o_param_abc.2638
"10101011110111100000000000000101",	-- 5446: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5447: 	lw	%ra, [%sp + 4]
"10010011110000000000000000000011",	-- 5448: 	lf	%f0, [%sp + 3]
"10010011110000010000000000000010",	-- 5449: 	lf	%f1, [%sp + 2]
"10010011110000100000000000000001",	-- 5450: 	lf	%f2, [%sp + 1]
"00111111111111100000000000000100",	-- 5451: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5452: 	addi	%sp, %sp, 5
"01011000000000000000010110111111",	-- 5453: 	jal	veciprod2.2600
"10101011110111100000000000000101",	-- 5454: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5455: 	lw	%ra, [%sp + 4]
"00111011110000010000000000000000",	-- 5456: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000100",	-- 5457: 	sf	%f0, [%sp + 4]
"00111111111111100000000000000101",	-- 5458: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5459: 	addi	%sp, %sp, 6
"01011000000000000000011001010110",	-- 5460: 	jal	o_isinvert.2628
"10101011110111100000000000000110",	-- 5461: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5462: 	lw	%ra, [%sp + 5]
"10010011110000000000000000000100",	-- 5463: 	lf	%f0, [%sp + 4]
"00111100001111100000000000000101",	-- 5464: 	sw	%r1, [%sp + 5]
"00111111111111100000000000000110",	-- 5465: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5466: 	addi	%sp, %sp, 7
"01011000000000000000010011011101",	-- 5467: 	jal	fisneg.2524
"10101011110111100000000000000111",	-- 5468: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5469: 	lw	%ra, [%sp + 6]
"10000100000000010001000000000000",	-- 5470: 	add	%r2, %r0, %r1
"00111011110000010000000000000101",	-- 5471: 	lw	%r1, [%sp + 5]
"00111111111111100000000000000110",	-- 5472: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5473: 	addi	%sp, %sp, 7
"01011000000000000000010011111000",	-- 5474: 	jal	xor.2565
"10101011110111100000000000000111",	-- 5475: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5476: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5477: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5478: 	bneq	%r1, %r2, bneq_else.9075
"11001100000000010000000000000001",	-- 5479: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5480: 	jr	%ra
	-- bneq_else.9075:
"11001100000000010000000000000000",	-- 5481: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5482: 	jr	%ra
	-- is_second_outside.2829:
"00111100001111100000000000000000",	-- 5483: 	sw	%r1, [%sp + 0]
"00111111111111100000000000000001",	-- 5484: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 5485: 	addi	%sp, %sp, 2
"01011000000000000000110001111010",	-- 5486: 	jal	quadratic.2737
"10101011110111100000000000000010",	-- 5487: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 5488: 	lw	%ra, [%sp + 1]
"00111011110000010000000000000000",	-- 5489: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000001",	-- 5490: 	sf	%f0, [%sp + 1]
"00111111111111100000000000000010",	-- 5491: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 5492: 	addi	%sp, %sp, 3
"01011000000000000000011001010010",	-- 5493: 	jal	o_form.2624
"10101011110111100000000000000011",	-- 5494: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 5495: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000011",	-- 5496: 	lli	%r2, 3
"00101000001000100000000000000110",	-- 5497: 	bneq	%r1, %r2, bneq_else.9076
"00010100000000000000000000000000",	-- 5498: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 5499: 	lhif	%f0, 1.000000
"10010011110000010000000000000001",	-- 5500: 	lf	%f1, [%sp + 1]
"11100100001000000000000000000000",	-- 5501: 	subf	%f0, %f1, %f0
"01010100000000000001010110000000",	-- 5502: 	j	bneq_cont.9077
	-- bneq_else.9076:
"10010011110000000000000000000001",	-- 5503: 	lf	%f0, [%sp + 1]
	-- bneq_cont.9077:
"00111011110000010000000000000000",	-- 5504: 	lw	%r1, [%sp + 0]
"10110000000111100000000000000010",	-- 5505: 	sf	%f0, [%sp + 2]
"00111111111111100000000000000011",	-- 5506: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 5507: 	addi	%sp, %sp, 4
"01011000000000000000011001010110",	-- 5508: 	jal	o_isinvert.2628
"10101011110111100000000000000100",	-- 5509: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 5510: 	lw	%ra, [%sp + 3]
"10010011110000000000000000000010",	-- 5511: 	lf	%f0, [%sp + 2]
"00111100001111100000000000000011",	-- 5512: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 5513: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5514: 	addi	%sp, %sp, 5
"01011000000000000000010011011101",	-- 5515: 	jal	fisneg.2524
"10101011110111100000000000000101",	-- 5516: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5517: 	lw	%ra, [%sp + 4]
"10000100000000010001000000000000",	-- 5518: 	add	%r2, %r0, %r1
"00111011110000010000000000000011",	-- 5519: 	lw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 5520: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5521: 	addi	%sp, %sp, 5
"01011000000000000000010011111000",	-- 5522: 	jal	xor.2565
"10101011110111100000000000000101",	-- 5523: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5524: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000000",	-- 5525: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5526: 	bneq	%r1, %r2, bneq_else.9078
"11001100000000010000000000000001",	-- 5527: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5528: 	jr	%ra
	-- bneq_else.9078:
"11001100000000010000000000000000",	-- 5529: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5530: 	jr	%ra
	-- is_outside.2834:
"10110000010111100000000000000000",	-- 5531: 	sf	%f2, [%sp + 0]
"10110000001111100000000000000001",	-- 5532: 	sf	%f1, [%sp + 1]
"00111100001111100000000000000010",	-- 5533: 	sw	%r1, [%sp + 2]
"10110000000111100000000000000011",	-- 5534: 	sf	%f0, [%sp + 3]
"00111111111111100000000000000100",	-- 5535: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 5536: 	addi	%sp, %sp, 5
"01011000000000000000011001101011",	-- 5537: 	jal	o_param_x.2640
"10101011110111100000000000000101",	-- 5538: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 5539: 	lw	%ra, [%sp + 4]
"10010011110000010000000000000011",	-- 5540: 	lf	%f1, [%sp + 3]
"11100100001000000000000000000000",	-- 5541: 	subf	%f0, %f1, %f0
"00111011110000010000000000000010",	-- 5542: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000100",	-- 5543: 	sf	%f0, [%sp + 4]
"00111111111111100000000000000101",	-- 5544: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 5545: 	addi	%sp, %sp, 6
"01011000000000000000011001110000",	-- 5546: 	jal	o_param_y.2642
"10101011110111100000000000000110",	-- 5547: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 5548: 	lw	%ra, [%sp + 5]
"10010011110000010000000000000001",	-- 5549: 	lf	%f1, [%sp + 1]
"11100100001000000000000000000000",	-- 5550: 	subf	%f0, %f1, %f0
"00111011110000010000000000000010",	-- 5551: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000101",	-- 5552: 	sf	%f0, [%sp + 5]
"00111111111111100000000000000110",	-- 5553: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5554: 	addi	%sp, %sp, 7
"01011000000000000000011001110101",	-- 5555: 	jal	o_param_z.2644
"10101011110111100000000000000111",	-- 5556: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5557: 	lw	%ra, [%sp + 6]
"10010011110000010000000000000000",	-- 5558: 	lf	%f1, [%sp + 0]
"11100100001000000000000000000000",	-- 5559: 	subf	%f0, %f1, %f0
"00111011110000010000000000000010",	-- 5560: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000110",	-- 5561: 	sf	%f0, [%sp + 6]
"00111111111111100000000000000111",	-- 5562: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 5563: 	addi	%sp, %sp, 8
"01011000000000000000011001010010",	-- 5564: 	jal	o_form.2624
"10101011110111100000000000001000",	-- 5565: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 5566: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000001",	-- 5567: 	lli	%r2, 1
"00101000001000100000000000000110",	-- 5568: 	bneq	%r1, %r2, bneq_else.9079
"10010011110000000000000000000100",	-- 5569: 	lf	%f0, [%sp + 4]
"10010011110000010000000000000101",	-- 5570: 	lf	%f1, [%sp + 5]
"10010011110000100000000000000110",	-- 5571: 	lf	%f2, [%sp + 6]
"00111011110000010000000000000010",	-- 5572: 	lw	%r1, [%sp + 2]
"01010100000000000001010011101001",	-- 5573: 	j	is_rect_outside.2819
	-- bneq_else.9079:
"11001100000000100000000000000010",	-- 5574: 	lli	%r2, 2
"00101000001000100000000000000110",	-- 5575: 	bneq	%r1, %r2, bneq_else.9080
"10010011110000000000000000000100",	-- 5576: 	lf	%f0, [%sp + 4]
"10010011110000010000000000000101",	-- 5577: 	lf	%f1, [%sp + 5]
"10010011110000100000000000000110",	-- 5578: 	lf	%f2, [%sp + 6]
"00111011110000010000000000000010",	-- 5579: 	lw	%r1, [%sp + 2]
"01010100000000000001010100111111",	-- 5580: 	j	is_plane_outside.2824
	-- bneq_else.9080:
"10010011110000000000000000000100",	-- 5581: 	lf	%f0, [%sp + 4]
"10010011110000010000000000000101",	-- 5582: 	lf	%f1, [%sp + 5]
"10010011110000100000000000000110",	-- 5583: 	lf	%f2, [%sp + 6]
"00111011110000010000000000000010",	-- 5584: 	lw	%r1, [%sp + 2]
"01010100000000000001010101101011",	-- 5585: 	j	is_second_outside.2829
	-- check_all_inside.2839:
"00111011011000110000000000000001",	-- 5586: 	lw	%r3, [%r27 + 1]
"10000100010000010010000000000000",	-- 5587: 	add	%r4, %r2, %r1
"00111000100001000000000000000000",	-- 5588: 	lw	%r4, [%r4 + 0]
"11001100000001011111111111111111",	-- 5589: 	lli	%r5, -1
"11001000000001011111111111111111",	-- 5590: 	lhi	%r5, -1
"00101000100001010000000000000011",	-- 5591: 	bneq	%r4, %r5, bneq_else.9081
"11001100000000010000000000000001",	-- 5592: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5593: 	jr	%ra
	-- bneq_else.9081:
"10000100011001000001100000000000",	-- 5594: 	add	%r3, %r3, %r4
"00111000011000110000000000000000",	-- 5595: 	lw	%r3, [%r3 + 0]
"10110000010111100000000000000000",	-- 5596: 	sf	%f2, [%sp + 0]
"10110000001111100000000000000001",	-- 5597: 	sf	%f1, [%sp + 1]
"10110000000111100000000000000010",	-- 5598: 	sf	%f0, [%sp + 2]
"00111100010111100000000000000011",	-- 5599: 	sw	%r2, [%sp + 3]
"00111111011111100000000000000100",	-- 5600: 	sw	%r27, [%sp + 4]
"00111100001111100000000000000101",	-- 5601: 	sw	%r1, [%sp + 5]
"10000100000000110000100000000000",	-- 5602: 	add	%r1, %r0, %r3
"00111111111111100000000000000110",	-- 5603: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5604: 	addi	%sp, %sp, 7
"01011000000000000001010110011011",	-- 5605: 	jal	is_outside.2834
"10101011110111100000000000000111",	-- 5606: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5607: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5608: 	lli	%r2, 0
"00101000001000100000000000001011",	-- 5609: 	bneq	%r1, %r2, bneq_else.9082
"11001100000000010000000000000001",	-- 5610: 	lli	%r1, 1
"00111011110000100000000000000101",	-- 5611: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 5612: 	add	%r1, %r2, %r1
"10010011110000000000000000000010",	-- 5613: 	lf	%f0, [%sp + 2]
"10010011110000010000000000000001",	-- 5614: 	lf	%f1, [%sp + 1]
"10010011110000100000000000000000",	-- 5615: 	lf	%f2, [%sp + 0]
"00111011110000100000000000000011",	-- 5616: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000100",	-- 5617: 	lw	%r27, [%sp + 4]
"00111011011110100000000000000000",	-- 5618: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5619: 	jr	%r26
	-- bneq_else.9082:
"11001100000000010000000000000000",	-- 5620: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5621: 	jr	%ra
	-- shadow_check_and_group.2845:
"00111011011000110000000000000111",	-- 5622: 	lw	%r3, [%r27 + 7]
"00111011011001000000000000000110",	-- 5623: 	lw	%r4, [%r27 + 6]
"00111011011001010000000000000101",	-- 5624: 	lw	%r5, [%r27 + 5]
"00111011011001100000000000000100",	-- 5625: 	lw	%r6, [%r27 + 4]
"00111011011001110000000000000011",	-- 5626: 	lw	%r7, [%r27 + 3]
"00111011011010000000000000000010",	-- 5627: 	lw	%r8, [%r27 + 2]
"00111011011010010000000000000001",	-- 5628: 	lw	%r9, [%r27 + 1]
"10000100010000010101000000000000",	-- 5629: 	add	%r10, %r2, %r1
"00111001010010100000000000000000",	-- 5630: 	lw	%r10, [%r10 + 0]
"11001100000010111111111111111111",	-- 5631: 	lli	%r11, -1
"11001000000010111111111111111111",	-- 5632: 	lhi	%r11, -1
"00101001010010110000000000000011",	-- 5633: 	bneq	%r10, %r11, bneq_else.9083
"11001100000000010000000000000000",	-- 5634: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5635: 	jr	%ra
	-- bneq_else.9083:
"10000100010000010101000000000000",	-- 5636: 	add	%r10, %r2, %r1
"00111001010010100000000000000000",	-- 5637: 	lw	%r10, [%r10 + 0]
"00111101001111100000000000000000",	-- 5638: 	sw	%r9, [%sp + 0]
"00111101000111100000000000000001",	-- 5639: 	sw	%r8, [%sp + 1]
"00111100111111100000000000000010",	-- 5640: 	sw	%r7, [%sp + 2]
"00111100010111100000000000000011",	-- 5641: 	sw	%r2, [%sp + 3]
"00111111011111100000000000000100",	-- 5642: 	sw	%r27, [%sp + 4]
"00111100001111100000000000000101",	-- 5643: 	sw	%r1, [%sp + 5]
"00111101010111100000000000000110",	-- 5644: 	sw	%r10, [%sp + 6]
"00111100101111100000000000000111",	-- 5645: 	sw	%r5, [%sp + 7]
"00111100100111100000000000001000",	-- 5646: 	sw	%r4, [%sp + 8]
"10000100000001100001000000000000",	-- 5647: 	add	%r2, %r0, %r6
"10000100000010100000100000000000",	-- 5648: 	add	%r1, %r0, %r10
"10000100000000111101100000000000",	-- 5649: 	add	%r27, %r0, %r3
"10000100000010000001100000000000",	-- 5650: 	add	%r3, %r0, %r8
"00111111111111100000000000001001",	-- 5651: 	sw	%ra, [%sp + 9]
"00111011011110100000000000000000",	-- 5652: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001010",	-- 5653: 	addi	%sp, %sp, 10
"01010011010000000000000000000000",	-- 5654: 	jalr	%r26
"10101011110111100000000000001010",	-- 5655: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 5656: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000000",	-- 5657: 	lli	%r2, 0
"00111011110000110000000000001000",	-- 5658: 	lw	%r3, [%sp + 8]
"10000100011000100001000000000000",	-- 5659: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 5660: 	lf	%f0, [%r2 + 0]
"11001100000000100000000000000000",	-- 5661: 	lli	%r2, 0
"10110000000111100000000000001001",	-- 5662: 	sf	%f0, [%sp + 9]
"00101000001000100000000000000011",	-- 5663: 	bneq	%r1, %r2, bneq_else.9084
"11001100000000010000000000000000",	-- 5664: 	lli	%r1, 0
"01010100000000000001011000101001",	-- 5665: 	j	bneq_cont.9085
	-- bneq_else.9084:
"00010100000000011100110011001101",	-- 5666: 	llif	%f1, -0.200000
"00010000000000011011111001001100",	-- 5667: 	lhif	%f1, -0.200000
"00111111111111100000000000001010",	-- 5668: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 5669: 	addi	%sp, %sp, 11
"01011000000000000000010011110011",	-- 5670: 	jal	fless.2532
"10101011110111100000000000001011",	-- 5671: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 5672: 	lw	%ra, [%sp + 10]
	-- bneq_cont.9085:
"11001100000000100000000000000000",	-- 5673: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 5674: 	bneq	%r1, %r2, bneq_else.9086
"00111011110000010000000000000110",	-- 5675: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000111",	-- 5676: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 5677: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 5678: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001010",	-- 5679: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 5680: 	addi	%sp, %sp, 11
"01011000000000000000011001010110",	-- 5681: 	jal	o_isinvert.2628
"10101011110111100000000000001011",	-- 5682: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 5683: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 5684: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5685: 	bneq	%r1, %r2, bneq_else.9087
"11001100000000010000000000000000",	-- 5686: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5687: 	jr	%ra
	-- bneq_else.9087:
"11001100000000010000000000000001",	-- 5688: 	lli	%r1, 1
"00111011110000100000000000000101",	-- 5689: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 5690: 	add	%r1, %r2, %r1
"00111011110000100000000000000011",	-- 5691: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000100",	-- 5692: 	lw	%r27, [%sp + 4]
"00111011011110100000000000000000",	-- 5693: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5694: 	jr	%r26
	-- bneq_else.9086:
"00010100000000001101011100001010",	-- 5695: 	llif	%f0, 0.010000
"00010000000000000011110000100011",	-- 5696: 	lhif	%f0, 0.010000
"10010011110000010000000000001001",	-- 5697: 	lf	%f1, [%sp + 9]
"11100000001000000000000000000000",	-- 5698: 	addf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 5699: 	lli	%r1, 0
"00111011110000100000000000000010",	-- 5700: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 5701: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 5702: 	lf	%f1, [%r1 + 0]
"11101000001000000000100000000000",	-- 5703: 	mulf	%f1, %f1, %f0
"11001100000000010000000000000000",	-- 5704: 	lli	%r1, 0
"00111011110000110000000000000001",	-- 5705: 	lw	%r3, [%sp + 1]
"10000100011000010000100000000000",	-- 5706: 	add	%r1, %r3, %r1
"10010000001000100000000000000000",	-- 5707: 	lf	%f2, [%r1 + 0]
"11100000001000100000100000000000",	-- 5708: 	addf	%f1, %f1, %f2
"11001100000000010000000000000001",	-- 5709: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 5710: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 5711: 	lf	%f2, [%r1 + 0]
"11101000010000000001000000000000",	-- 5712: 	mulf	%f2, %f2, %f0
"11001100000000010000000000000001",	-- 5713: 	lli	%r1, 1
"10000100011000010000100000000000",	-- 5714: 	add	%r1, %r3, %r1
"10010000001000110000000000000000",	-- 5715: 	lf	%f3, [%r1 + 0]
"11100000010000110001000000000000",	-- 5716: 	addf	%f2, %f2, %f3
"11001100000000010000000000000010",	-- 5717: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 5718: 	add	%r1, %r2, %r1
"10010000001000110000000000000000",	-- 5719: 	lf	%f3, [%r1 + 0]
"11101000011000000000000000000000",	-- 5720: 	mulf	%f0, %f3, %f0
"11001100000000010000000000000010",	-- 5721: 	lli	%r1, 2
"10000100011000010000100000000000",	-- 5722: 	add	%r1, %r3, %r1
"10010000001000110000000000000000",	-- 5723: 	lf	%f3, [%r1 + 0]
"11100000000000110000000000000000",	-- 5724: 	addf	%f0, %f0, %f3
"11001100000000010000000000000000",	-- 5725: 	lli	%r1, 0
"00111011110000100000000000000011",	-- 5726: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000000",	-- 5727: 	lw	%r27, [%sp + 0]
"00001100010111110000000000000000",	-- 5728: 	movf	%f31, %f2
"00001100000000100000000000000000",	-- 5729: 	movf	%f2, %f0
"00001100001000000000000000000000",	-- 5730: 	movf	%f0, %f1
"00001111111000010000000000000000",	-- 5731: 	movf	%f1, %f31
"00111111111111100000000000001010",	-- 5732: 	sw	%ra, [%sp + 10]
"00111011011110100000000000000000",	-- 5733: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001011",	-- 5734: 	addi	%sp, %sp, 11
"01010011010000000000000000000000",	-- 5735: 	jalr	%r26
"10101011110111100000000000001011",	-- 5736: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 5737: 	lw	%ra, [%sp + 10]
"11001100000000100000000000000000",	-- 5738: 	lli	%r2, 0
"00101000001000100000000000001000",	-- 5739: 	bneq	%r1, %r2, bneq_else.9088
"11001100000000010000000000000001",	-- 5740: 	lli	%r1, 1
"00111011110000100000000000000101",	-- 5741: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 5742: 	add	%r1, %r2, %r1
"00111011110000100000000000000011",	-- 5743: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000100",	-- 5744: 	lw	%r27, [%sp + 4]
"00111011011110100000000000000000",	-- 5745: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5746: 	jr	%r26
	-- bneq_else.9088:
"11001100000000010000000000000001",	-- 5747: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5748: 	jr	%ra
	-- shadow_check_one_or_group.2848:
"00111011011000110000000000000010",	-- 5749: 	lw	%r3, [%r27 + 2]
"00111011011001000000000000000001",	-- 5750: 	lw	%r4, [%r27 + 1]
"10000100010000010010100000000000",	-- 5751: 	add	%r5, %r2, %r1
"00111000101001010000000000000000",	-- 5752: 	lw	%r5, [%r5 + 0]
"11001100000001101111111111111111",	-- 5753: 	lli	%r6, -1
"11001000000001101111111111111111",	-- 5754: 	lhi	%r6, -1
"00101000101001100000000000000011",	-- 5755: 	bneq	%r5, %r6, bneq_else.9089
"11001100000000010000000000000000",	-- 5756: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5757: 	jr	%ra
	-- bneq_else.9089:
"10000100100001010010000000000000",	-- 5758: 	add	%r4, %r4, %r5
"00111000100001000000000000000000",	-- 5759: 	lw	%r4, [%r4 + 0]
"11001100000001010000000000000000",	-- 5760: 	lli	%r5, 0
"00111100010111100000000000000000",	-- 5761: 	sw	%r2, [%sp + 0]
"00111111011111100000000000000001",	-- 5762: 	sw	%r27, [%sp + 1]
"00111100001111100000000000000010",	-- 5763: 	sw	%r1, [%sp + 2]
"10000100000001000001000000000000",	-- 5764: 	add	%r2, %r0, %r4
"10000100000001010000100000000000",	-- 5765: 	add	%r1, %r0, %r5
"10000100000000111101100000000000",	-- 5766: 	add	%r27, %r0, %r3
"00111111111111100000000000000011",	-- 5767: 	sw	%ra, [%sp + 3]
"00111011011110100000000000000000",	-- 5768: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000100",	-- 5769: 	addi	%sp, %sp, 4
"01010011010000000000000000000000",	-- 5770: 	jalr	%r26
"10101011110111100000000000000100",	-- 5771: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 5772: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000000",	-- 5773: 	lli	%r2, 0
"00101000001000100000000000001000",	-- 5774: 	bneq	%r1, %r2, bneq_else.9090
"11001100000000010000000000000001",	-- 5775: 	lli	%r1, 1
"00111011110000100000000000000010",	-- 5776: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 5777: 	add	%r1, %r2, %r1
"00111011110000100000000000000000",	-- 5778: 	lw	%r2, [%sp + 0]
"00111011110110110000000000000001",	-- 5779: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 5780: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5781: 	jr	%r26
	-- bneq_else.9090:
"11001100000000010000000000000001",	-- 5782: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5783: 	jr	%ra
	-- shadow_check_one_or_matrix.2851:
"00111011011000110000000000000101",	-- 5784: 	lw	%r3, [%r27 + 5]
"00111011011001000000000000000100",	-- 5785: 	lw	%r4, [%r27 + 4]
"00111011011001010000000000000011",	-- 5786: 	lw	%r5, [%r27 + 3]
"00111011011001100000000000000010",	-- 5787: 	lw	%r6, [%r27 + 2]
"00111011011001110000000000000001",	-- 5788: 	lw	%r7, [%r27 + 1]
"10000100010000010100000000000000",	-- 5789: 	add	%r8, %r2, %r1
"00111001000010000000000000000000",	-- 5790: 	lw	%r8, [%r8 + 0]
"11001100000010010000000000000000",	-- 5791: 	lli	%r9, 0
"10000101000010010100100000000000",	-- 5792: 	add	%r9, %r8, %r9
"00111001001010010000000000000000",	-- 5793: 	lw	%r9, [%r9 + 0]
"11001100000010101111111111111111",	-- 5794: 	lli	%r10, -1
"11001000000010101111111111111111",	-- 5795: 	lhi	%r10, -1
"00101001001010100000000000000011",	-- 5796: 	bneq	%r9, %r10, bneq_else.9091
"11001100000000010000000000000000",	-- 5797: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 5798: 	jr	%ra
	-- bneq_else.9091:
"11001100000010100000000001100011",	-- 5799: 	lli	%r10, 99
"00111101000111100000000000000000",	-- 5800: 	sw	%r8, [%sp + 0]
"00111100101111100000000000000001",	-- 5801: 	sw	%r5, [%sp + 1]
"00111100010111100000000000000010",	-- 5802: 	sw	%r2, [%sp + 2]
"00111111011111100000000000000011",	-- 5803: 	sw	%r27, [%sp + 3]
"00111100001111100000000000000100",	-- 5804: 	sw	%r1, [%sp + 4]
"00101001001010100000000000000011",	-- 5805: 	bneq	%r9, %r10, bneq_else.9092
"11001100000000010000000000000001",	-- 5806: 	lli	%r1, 1
"01010100000000000001011011011100",	-- 5807: 	j	bneq_cont.9093
	-- bneq_else.9092:
"00111100100111100000000000000101",	-- 5808: 	sw	%r4, [%sp + 5]
"10000100000001100001000000000000",	-- 5809: 	add	%r2, %r0, %r6
"10000100000010010000100000000000",	-- 5810: 	add	%r1, %r0, %r9
"10000100000000111101100000000000",	-- 5811: 	add	%r27, %r0, %r3
"10000100000001110001100000000000",	-- 5812: 	add	%r3, %r0, %r7
"00111111111111100000000000000110",	-- 5813: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 5814: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 5815: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 5816: 	jalr	%r26
"10101011110111100000000000000111",	-- 5817: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5818: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5819: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5820: 	bneq	%r1, %r2, bneq_else.9094
"11001100000000010000000000000000",	-- 5821: 	lli	%r1, 0
"01010100000000000001011011011100",	-- 5822: 	j	bneq_cont.9095
	-- bneq_else.9094:
"11001100000000010000000000000000",	-- 5823: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 5824: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 5825: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 5826: 	lf	%f0, [%r1 + 0]
"00010100000000011100110011001101",	-- 5827: 	llif	%f1, -0.100000
"00010000000000011011110111001100",	-- 5828: 	lhif	%f1, -0.100000
"00111111111111100000000000000110",	-- 5829: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 5830: 	addi	%sp, %sp, 7
"01011000000000000000010011110011",	-- 5831: 	jal	fless.2532
"10101011110111100000000000000111",	-- 5832: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5833: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5834: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5835: 	bneq	%r1, %r2, bneq_else.9096
"11001100000000010000000000000000",	-- 5836: 	lli	%r1, 0
"01010100000000000001011011011100",	-- 5837: 	j	bneq_cont.9097
	-- bneq_else.9096:
"11001100000000010000000000000001",	-- 5838: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 5839: 	lw	%r2, [%sp + 0]
"00111011110110110000000000000001",	-- 5840: 	lw	%r27, [%sp + 1]
"00111111111111100000000000000110",	-- 5841: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 5842: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 5843: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 5844: 	jalr	%r26
"10101011110111100000000000000111",	-- 5845: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5846: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5847: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 5848: 	bneq	%r1, %r2, bneq_else.9098
"11001100000000010000000000000000",	-- 5849: 	lli	%r1, 0
"01010100000000000001011011011100",	-- 5850: 	j	bneq_cont.9099
	-- bneq_else.9098:
"11001100000000010000000000000001",	-- 5851: 	lli	%r1, 1
	-- bneq_cont.9099:
	-- bneq_cont.9097:
	-- bneq_cont.9095:
	-- bneq_cont.9093:
"11001100000000100000000000000000",	-- 5852: 	lli	%r2, 0
"00101000001000100000000000001000",	-- 5853: 	bneq	%r1, %r2, bneq_else.9100
"11001100000000010000000000000001",	-- 5854: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 5855: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5856: 	add	%r1, %r2, %r1
"00111011110000100000000000000010",	-- 5857: 	lw	%r2, [%sp + 2]
"00111011110110110000000000000011",	-- 5858: 	lw	%r27, [%sp + 3]
"00111011011110100000000000000000",	-- 5859: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5860: 	jr	%r26
	-- bneq_else.9100:
"11001100000000010000000000000001",	-- 5861: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 5862: 	lw	%r2, [%sp + 0]
"00111011110110110000000000000001",	-- 5863: 	lw	%r27, [%sp + 1]
"00111111111111100000000000000110",	-- 5864: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 5865: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 5866: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 5867: 	jalr	%r26
"10101011110111100000000000000111",	-- 5868: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 5869: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 5870: 	lli	%r2, 0
"00101000001000100000000000001000",	-- 5871: 	bneq	%r1, %r2, bneq_else.9101
"11001100000000010000000000000001",	-- 5872: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 5873: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 5874: 	add	%r1, %r2, %r1
"00111011110000100000000000000010",	-- 5875: 	lw	%r2, [%sp + 2]
"00111011110110110000000000000011",	-- 5876: 	lw	%r27, [%sp + 3]
"00111011011110100000000000000000",	-- 5877: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5878: 	jr	%r26
	-- bneq_else.9101:
"11001100000000010000000000000001",	-- 5879: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 5880: 	jr	%ra
	-- solve_each_element.2854:
"00111011011001000000000000001001",	-- 5881: 	lw	%r4, [%r27 + 9]
"00111011011001010000000000001000",	-- 5882: 	lw	%r5, [%r27 + 8]
"00111011011001100000000000000111",	-- 5883: 	lw	%r6, [%r27 + 7]
"00111011011001110000000000000110",	-- 5884: 	lw	%r7, [%r27 + 6]
"00111011011010000000000000000101",	-- 5885: 	lw	%r8, [%r27 + 5]
"00111011011010010000000000000100",	-- 5886: 	lw	%r9, [%r27 + 4]
"00111011011010100000000000000011",	-- 5887: 	lw	%r10, [%r27 + 3]
"00111011011010110000000000000010",	-- 5888: 	lw	%r11, [%r27 + 2]
"00111011011011000000000000000001",	-- 5889: 	lw	%r12, [%r27 + 1]
"10000100010000010110100000000000",	-- 5890: 	add	%r13, %r2, %r1
"00111001101011010000000000000000",	-- 5891: 	lw	%r13, [%r13 + 0]
"11001100000011101111111111111111",	-- 5892: 	lli	%r14, -1
"11001000000011101111111111111111",	-- 5893: 	lhi	%r14, -1
"00101001101011100000000000000010",	-- 5894: 	bneq	%r13, %r14, bneq_else.9102
"01001111111000000000000000000000",	-- 5895: 	jr	%ra
	-- bneq_else.9102:
"00111101001111100000000000000000",	-- 5896: 	sw	%r9, [%sp + 0]
"00111101011111100000000000000001",	-- 5897: 	sw	%r11, [%sp + 1]
"00111101010111100000000000000010",	-- 5898: 	sw	%r10, [%sp + 2]
"00111101100111100000000000000011",	-- 5899: 	sw	%r12, [%sp + 3]
"00111100101111100000000000000100",	-- 5900: 	sw	%r5, [%sp + 4]
"00111100100111100000000000000101",	-- 5901: 	sw	%r4, [%sp + 5]
"00111100110111100000000000000110",	-- 5902: 	sw	%r6, [%sp + 6]
"00111100011111100000000000000111",	-- 5903: 	sw	%r3, [%sp + 7]
"00111100010111100000000000001000",	-- 5904: 	sw	%r2, [%sp + 8]
"00111111011111100000000000001001",	-- 5905: 	sw	%r27, [%sp + 9]
"00111100001111100000000000001010",	-- 5906: 	sw	%r1, [%sp + 10]
"00111101101111100000000000001011",	-- 5907: 	sw	%r13, [%sp + 11]
"00111101000111100000000000001100",	-- 5908: 	sw	%r8, [%sp + 12]
"10000100000000110001000000000000",	-- 5909: 	add	%r2, %r0, %r3
"10000100000011010000100000000000",	-- 5910: 	add	%r1, %r0, %r13
"10000100000001111101100000000000",	-- 5911: 	add	%r27, %r0, %r7
"10000100000001010001100000000000",	-- 5912: 	add	%r3, %r0, %r5
"00111111111111100000000000001101",	-- 5913: 	sw	%ra, [%sp + 13]
"00111011011110100000000000000000",	-- 5914: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001110",	-- 5915: 	addi	%sp, %sp, 14
"01010011010000000000000000000000",	-- 5916: 	jalr	%r26
"10101011110111100000000000001110",	-- 5917: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 5918: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 5919: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 5920: 	bneq	%r1, %r2, bneq_else.9104
"00111011110000010000000000001011",	-- 5921: 	lw	%r1, [%sp + 11]
"00111011110000100000000000001100",	-- 5922: 	lw	%r2, [%sp + 12]
"10000100010000010000100000000000",	-- 5923: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 5924: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001101",	-- 5925: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 5926: 	addi	%sp, %sp, 14
"01011000000000000000011001010110",	-- 5927: 	jal	o_isinvert.2628
"10101011110111100000000000001110",	-- 5928: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 5929: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 5930: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 5931: 	bneq	%r1, %r2, bneq_else.9105
"01001111111000000000000000000000",	-- 5932: 	jr	%ra
	-- bneq_else.9105:
"11001100000000010000000000000001",	-- 5933: 	lli	%r1, 1
"00111011110000100000000000001010",	-- 5934: 	lw	%r2, [%sp + 10]
"10000100010000010000100000000000",	-- 5935: 	add	%r1, %r2, %r1
"00111011110000100000000000001000",	-- 5936: 	lw	%r2, [%sp + 8]
"00111011110000110000000000000111",	-- 5937: 	lw	%r3, [%sp + 7]
"00111011110110110000000000001001",	-- 5938: 	lw	%r27, [%sp + 9]
"00111011011110100000000000000000",	-- 5939: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 5940: 	jr	%r26
	-- bneq_else.9104:
"11001100000000100000000000000000",	-- 5941: 	lli	%r2, 0
"00111011110000110000000000000110",	-- 5942: 	lw	%r3, [%sp + 6]
"10000100011000100001000000000000",	-- 5943: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 5944: 	lf	%f1, [%r2 + 0]
"00010100000000000000000000000000",	-- 5945: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 5946: 	lhif	%f0, 0.000000
"00111100001111100000000000001101",	-- 5947: 	sw	%r1, [%sp + 13]
"10110000001111100000000000001110",	-- 5948: 	sf	%f1, [%sp + 14]
"00111111111111100000000000001111",	-- 5949: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 5950: 	addi	%sp, %sp, 16
"01011000000000000000010011110011",	-- 5951: 	jal	fless.2532
"10101011110111100000000000010000",	-- 5952: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 5953: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 5954: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 5955: 	bneq	%r1, %r2, bneq_else.9107
"01010100000000000001011110011100",	-- 5956: 	j	bneq_cont.9108
	-- bneq_else.9107:
"11001100000000010000000000000000",	-- 5957: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 5958: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 5959: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 5960: 	lf	%f1, [%r1 + 0]
"10010011110000000000000000001110",	-- 5961: 	lf	%f0, [%sp + 14]
"00111111111111100000000000001111",	-- 5962: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 5963: 	addi	%sp, %sp, 16
"01011000000000000000010011110011",	-- 5964: 	jal	fless.2532
"10101011110111100000000000010000",	-- 5965: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 5966: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 5967: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 5968: 	bneq	%r1, %r2, bneq_else.9109
"01010100000000000001011110011100",	-- 5969: 	j	bneq_cont.9110
	-- bneq_else.9109:
"00010100000000001101011100001010",	-- 5970: 	llif	%f0, 0.010000
"00010000000000000011110000100011",	-- 5971: 	lhif	%f0, 0.010000
"10010011110000010000000000001110",	-- 5972: 	lf	%f1, [%sp + 14]
"11100000001000000000000000000000",	-- 5973: 	addf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 5974: 	lli	%r1, 0
"00111011110000100000000000000111",	-- 5975: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 5976: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 5977: 	lf	%f1, [%r1 + 0]
"11101000001000000000100000000000",	-- 5978: 	mulf	%f1, %f1, %f0
"11001100000000010000000000000000",	-- 5979: 	lli	%r1, 0
"00111011110000110000000000000100",	-- 5980: 	lw	%r3, [%sp + 4]
"10000100011000010000100000000000",	-- 5981: 	add	%r1, %r3, %r1
"10010000001000100000000000000000",	-- 5982: 	lf	%f2, [%r1 + 0]
"11100000001000100000100000000000",	-- 5983: 	addf	%f1, %f1, %f2
"11001100000000010000000000000001",	-- 5984: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 5985: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 5986: 	lf	%f2, [%r1 + 0]
"11101000010000000001000000000000",	-- 5987: 	mulf	%f2, %f2, %f0
"11001100000000010000000000000001",	-- 5988: 	lli	%r1, 1
"10000100011000010000100000000000",	-- 5989: 	add	%r1, %r3, %r1
"10010000001000110000000000000000",	-- 5990: 	lf	%f3, [%r1 + 0]
"11100000010000110001000000000000",	-- 5991: 	addf	%f2, %f2, %f3
"11001100000000010000000000000010",	-- 5992: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 5993: 	add	%r1, %r2, %r1
"10010000001000110000000000000000",	-- 5994: 	lf	%f3, [%r1 + 0]
"11101000011000000001100000000000",	-- 5995: 	mulf	%f3, %f3, %f0
"11001100000000010000000000000010",	-- 5996: 	lli	%r1, 2
"10000100011000010000100000000000",	-- 5997: 	add	%r1, %r3, %r1
"10010000001001000000000000000000",	-- 5998: 	lf	%f4, [%r1 + 0]
"11100000011001000001100000000000",	-- 5999: 	addf	%f3, %f3, %f4
"11001100000000010000000000000000",	-- 6000: 	lli	%r1, 0
"00111011110000110000000000001000",	-- 6001: 	lw	%r3, [%sp + 8]
"00111011110110110000000000000011",	-- 6002: 	lw	%r27, [%sp + 3]
"10110000011111100000000000001111",	-- 6003: 	sf	%f3, [%sp + 15]
"10110000010111100000000000010000",	-- 6004: 	sf	%f2, [%sp + 16]
"10110000001111100000000000010001",	-- 6005: 	sf	%f1, [%sp + 17]
"10110000000111100000000000010010",	-- 6006: 	sf	%f0, [%sp + 18]
"10000100000000110001000000000000",	-- 6007: 	add	%r2, %r0, %r3
"00001100001000000000000000000000",	-- 6008: 	movf	%f0, %f1
"00001100010000010000000000000000",	-- 6009: 	movf	%f1, %f2
"00001100011000100000000000000000",	-- 6010: 	movf	%f2, %f3
"00111111111111100000000000010011",	-- 6011: 	sw	%ra, [%sp + 19]
"00111011011110100000000000000000",	-- 6012: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010100",	-- 6013: 	addi	%sp, %sp, 20
"01010011010000000000000000000000",	-- 6014: 	jalr	%r26
"10101011110111100000000000010100",	-- 6015: 	subi	%sp, %sp, 20
"00111011110111110000000000010011",	-- 6016: 	lw	%ra, [%sp + 19]
"11001100000000100000000000000000",	-- 6017: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6018: 	bneq	%r1, %r2, bneq_else.9111
"01010100000000000001011110011100",	-- 6019: 	j	bneq_cont.9112
	-- bneq_else.9111:
"11001100000000010000000000000000",	-- 6020: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 6021: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 6022: 	add	%r1, %r2, %r1
"10010011110000000000000000010010",	-- 6023: 	lf	%f0, [%sp + 18]
"10110000000000010000000000000000",	-- 6024: 	sf	%f0, [%r1 + 0]
"10010011110000000000000000010001",	-- 6025: 	lf	%f0, [%sp + 17]
"10010011110000010000000000010000",	-- 6026: 	lf	%f1, [%sp + 16]
"10010011110000100000000000001111",	-- 6027: 	lf	%f2, [%sp + 15]
"00111011110000010000000000000010",	-- 6028: 	lw	%r1, [%sp + 2]
"00111111111111100000000000010011",	-- 6029: 	sw	%ra, [%sp + 19]
"10100111110111100000000000010100",	-- 6030: 	addi	%sp, %sp, 20
"01011000000000000000010100100110",	-- 6031: 	jal	vecset.2576
"10101011110111100000000000010100",	-- 6032: 	subi	%sp, %sp, 20
"00111011110111110000000000010011",	-- 6033: 	lw	%ra, [%sp + 19]
"11001100000000010000000000000000",	-- 6034: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 6035: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 6036: 	add	%r1, %r2, %r1
"00111011110000100000000000001011",	-- 6037: 	lw	%r2, [%sp + 11]
"00111100010000010000000000000000",	-- 6038: 	sw	%r2, [%r1 + 0]
"11001100000000010000000000000000",	-- 6039: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 6040: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6041: 	add	%r1, %r2, %r1
"00111011110000100000000000001101",	-- 6042: 	lw	%r2, [%sp + 13]
"00111100010000010000000000000000",	-- 6043: 	sw	%r2, [%r1 + 0]
	-- bneq_cont.9112:
	-- bneq_cont.9110:
	-- bneq_cont.9108:
"11001100000000010000000000000001",	-- 6044: 	lli	%r1, 1
"00111011110000100000000000001010",	-- 6045: 	lw	%r2, [%sp + 10]
"10000100010000010000100000000000",	-- 6046: 	add	%r1, %r2, %r1
"00111011110000100000000000001000",	-- 6047: 	lw	%r2, [%sp + 8]
"00111011110000110000000000000111",	-- 6048: 	lw	%r3, [%sp + 7]
"00111011110110110000000000001001",	-- 6049: 	lw	%r27, [%sp + 9]
"00111011011110100000000000000000",	-- 6050: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6051: 	jr	%r26
	-- solve_one_or_network.2858:
"00111011011001000000000000000010",	-- 6052: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 6053: 	lw	%r5, [%r27 + 1]
"10000100010000010011000000000000",	-- 6054: 	add	%r6, %r2, %r1
"00111000110001100000000000000000",	-- 6055: 	lw	%r6, [%r6 + 0]
"11001100000001111111111111111111",	-- 6056: 	lli	%r7, -1
"11001000000001111111111111111111",	-- 6057: 	lhi	%r7, -1
"00101000110001110000000000000010",	-- 6058: 	bneq	%r6, %r7, bneq_else.9113
"01001111111000000000000000000000",	-- 6059: 	jr	%ra
	-- bneq_else.9113:
"10000100101001100010100000000000",	-- 6060: 	add	%r5, %r5, %r6
"00111000101001010000000000000000",	-- 6061: 	lw	%r5, [%r5 + 0]
"11001100000001100000000000000000",	-- 6062: 	lli	%r6, 0
"00111100011111100000000000000000",	-- 6063: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 6064: 	sw	%r2, [%sp + 1]
"00111111011111100000000000000010",	-- 6065: 	sw	%r27, [%sp + 2]
"00111100001111100000000000000011",	-- 6066: 	sw	%r1, [%sp + 3]
"10000100000001010001000000000000",	-- 6067: 	add	%r2, %r0, %r5
"10000100000001100000100000000000",	-- 6068: 	add	%r1, %r0, %r6
"10000100000001001101100000000000",	-- 6069: 	add	%r27, %r0, %r4
"00111111111111100000000000000100",	-- 6070: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 6071: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 6072: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 6073: 	jalr	%r26
"10101011110111100000000000000101",	-- 6074: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6075: 	lw	%ra, [%sp + 4]
"11001100000000010000000000000001",	-- 6076: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 6077: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 6078: 	add	%r1, %r2, %r1
"00111011110000100000000000000001",	-- 6079: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 6080: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000010",	-- 6081: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 6082: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6083: 	jr	%r26
	-- trace_or_matrix.2862:
"00111011011001000000000000000101",	-- 6084: 	lw	%r4, [%r27 + 5]
"00111011011001010000000000000100",	-- 6085: 	lw	%r5, [%r27 + 4]
"00111011011001100000000000000011",	-- 6086: 	lw	%r6, [%r27 + 3]
"00111011011001110000000000000010",	-- 6087: 	lw	%r7, [%r27 + 2]
"00111011011010000000000000000001",	-- 6088: 	lw	%r8, [%r27 + 1]
"10000100010000010100100000000000",	-- 6089: 	add	%r9, %r2, %r1
"00111001001010010000000000000000",	-- 6090: 	lw	%r9, [%r9 + 0]
"11001100000010100000000000000000",	-- 6091: 	lli	%r10, 0
"10000101001010100101000000000000",	-- 6092: 	add	%r10, %r9, %r10
"00111001010010100000000000000000",	-- 6093: 	lw	%r10, [%r10 + 0]
"11001100000010111111111111111111",	-- 6094: 	lli	%r11, -1
"11001000000010111111111111111111",	-- 6095: 	lhi	%r11, -1
"00101001010010110000000000000010",	-- 6096: 	bneq	%r10, %r11, bneq_else.9115
"01001111111000000000000000000000",	-- 6097: 	jr	%ra
	-- bneq_else.9115:
"11001100000010110000000001100011",	-- 6098: 	lli	%r11, 99
"00111100011111100000000000000000",	-- 6099: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 6100: 	sw	%r2, [%sp + 1]
"00111111011111100000000000000010",	-- 6101: 	sw	%r27, [%sp + 2]
"00111100001111100000000000000011",	-- 6102: 	sw	%r1, [%sp + 3]
"00101001010010110000000000001100",	-- 6103: 	bneq	%r10, %r11, bneq_else.9117
"11001100000001000000000000000001",	-- 6104: 	lli	%r4, 1
"10000100000010010001000000000000",	-- 6105: 	add	%r2, %r0, %r9
"10000100000001000000100000000000",	-- 6106: 	add	%r1, %r0, %r4
"10000100000010001101100000000000",	-- 6107: 	add	%r27, %r0, %r8
"00111111111111100000000000000100",	-- 6108: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 6109: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 6110: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 6111: 	jalr	%r26
"10101011110111100000000000000101",	-- 6112: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6113: 	lw	%ra, [%sp + 4]
"01010100000000000001100000001110",	-- 6114: 	j	bneq_cont.9118
	-- bneq_else.9117:
"00111101001111100000000000000100",	-- 6115: 	sw	%r9, [%sp + 4]
"00111101000111100000000000000101",	-- 6116: 	sw	%r8, [%sp + 5]
"00111100100111100000000000000110",	-- 6117: 	sw	%r4, [%sp + 6]
"00111100110111100000000000000111",	-- 6118: 	sw	%r6, [%sp + 7]
"10000100000000110001000000000000",	-- 6119: 	add	%r2, %r0, %r3
"10000100000010100000100000000000",	-- 6120: 	add	%r1, %r0, %r10
"10000100000001111101100000000000",	-- 6121: 	add	%r27, %r0, %r7
"10000100000001010001100000000000",	-- 6122: 	add	%r3, %r0, %r5
"00111111111111100000000000001000",	-- 6123: 	sw	%ra, [%sp + 8]
"00111011011110100000000000000000",	-- 6124: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001001",	-- 6125: 	addi	%sp, %sp, 9
"01010011010000000000000000000000",	-- 6126: 	jalr	%r26
"10101011110111100000000000001001",	-- 6127: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6128: 	lw	%ra, [%sp + 8]
"11001100000000100000000000000000",	-- 6129: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6130: 	bneq	%r1, %r2, bneq_else.9119
"01010100000000000001100000001110",	-- 6131: 	j	bneq_cont.9120
	-- bneq_else.9119:
"11001100000000010000000000000000",	-- 6132: 	lli	%r1, 0
"00111011110000100000000000000111",	-- 6133: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 6134: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 6135: 	lf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 6136: 	lli	%r1, 0
"00111011110000100000000000000110",	-- 6137: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 6138: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6139: 	lf	%f1, [%r1 + 0]
"00111111111111100000000000001000",	-- 6140: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 6141: 	addi	%sp, %sp, 9
"01011000000000000000010011110011",	-- 6142: 	jal	fless.2532
"10101011110111100000000000001001",	-- 6143: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6144: 	lw	%ra, [%sp + 8]
"11001100000000100000000000000000",	-- 6145: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6146: 	bneq	%r1, %r2, bneq_else.9121
"01010100000000000001100000001110",	-- 6147: 	j	bneq_cont.9122
	-- bneq_else.9121:
"11001100000000010000000000000001",	-- 6148: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 6149: 	lw	%r2, [%sp + 4]
"00111011110000110000000000000000",	-- 6150: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000101",	-- 6151: 	lw	%r27, [%sp + 5]
"00111111111111100000000000001000",	-- 6152: 	sw	%ra, [%sp + 8]
"00111011011110100000000000000000",	-- 6153: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001001",	-- 6154: 	addi	%sp, %sp, 9
"01010011010000000000000000000000",	-- 6155: 	jalr	%r26
"10101011110111100000000000001001",	-- 6156: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6157: 	lw	%ra, [%sp + 8]
	-- bneq_cont.9122:
	-- bneq_cont.9120:
	-- bneq_cont.9118:
"11001100000000010000000000000001",	-- 6158: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 6159: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 6160: 	add	%r1, %r2, %r1
"00111011110000100000000000000001",	-- 6161: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 6162: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000010",	-- 6163: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 6164: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6165: 	jr	%r26
	-- judge_intersection.2866:
"00111011011000100000000000000011",	-- 6166: 	lw	%r2, [%r27 + 3]
"00111011011000110000000000000010",	-- 6167: 	lw	%r3, [%r27 + 2]
"00111011011001000000000000000001",	-- 6168: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 6169: 	lli	%r5, 0
"00010100000000000110101100101000",	-- 6170: 	llif	%f0, 1000000000.000000
"00010000000000000100111001101110",	-- 6171: 	lhif	%f0, 1000000000.000000
"10000100011001010010100000000000",	-- 6172: 	add	%r5, %r3, %r5
"10110000000001010000000000000000",	-- 6173: 	sf	%f0, [%r5 + 0]
"11001100000001010000000000000000",	-- 6174: 	lli	%r5, 0
"11001100000001100000000000000000",	-- 6175: 	lli	%r6, 0
"10000100100001100010000000000000",	-- 6176: 	add	%r4, %r4, %r6
"00111000100001000000000000000000",	-- 6177: 	lw	%r4, [%r4 + 0]
"00111100011111100000000000000000",	-- 6178: 	sw	%r3, [%sp + 0]
"10000100000000010001100000000000",	-- 6179: 	add	%r3, %r0, %r1
"10000100000000101101100000000000",	-- 6180: 	add	%r27, %r0, %r2
"10000100000001000001000000000000",	-- 6181: 	add	%r2, %r0, %r4
"10000100000001010000100000000000",	-- 6182: 	add	%r1, %r0, %r5
"00111111111111100000000000000001",	-- 6183: 	sw	%ra, [%sp + 1]
"00111011011110100000000000000000",	-- 6184: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000010",	-- 6185: 	addi	%sp, %sp, 2
"01010011010000000000000000000000",	-- 6186: 	jalr	%r26
"10101011110111100000000000000010",	-- 6187: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 6188: 	lw	%ra, [%sp + 1]
"11001100000000010000000000000000",	-- 6189: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 6190: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6191: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6192: 	lf	%f1, [%r1 + 0]
"00010100000000001100110011001101",	-- 6193: 	llif	%f0, -0.100000
"00010000000000001011110111001100",	-- 6194: 	lhif	%f0, -0.100000
"10110000001111100000000000000001",	-- 6195: 	sf	%f1, [%sp + 1]
"00111111111111100000000000000010",	-- 6196: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 6197: 	addi	%sp, %sp, 3
"01011000000000000000010011110011",	-- 6198: 	jal	fless.2532
"10101011110111100000000000000011",	-- 6199: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 6200: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000000",	-- 6201: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 6202: 	bneq	%r1, %r2, bneq_else.9123
"11001100000000010000000000000000",	-- 6203: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 6204: 	jr	%ra
	-- bneq_else.9123:
"00010100000000011011110000100000",	-- 6205: 	llif	%f1, 100000000.000000
"00010000000000010100110010111110",	-- 6206: 	lhif	%f1, 100000000.000000
"10010011110000000000000000000001",	-- 6207: 	lf	%f0, [%sp + 1]
"01010100000000000000010011110011",	-- 6208: 	j	fless.2532
	-- solve_each_element_fast.2868:
"00111011011001000000000000001001",	-- 6209: 	lw	%r4, [%r27 + 9]
"00111011011001010000000000001000",	-- 6210: 	lw	%r5, [%r27 + 8]
"00111011011001100000000000000111",	-- 6211: 	lw	%r6, [%r27 + 7]
"00111011011001110000000000000110",	-- 6212: 	lw	%r7, [%r27 + 6]
"00111011011010000000000000000101",	-- 6213: 	lw	%r8, [%r27 + 5]
"00111011011010010000000000000100",	-- 6214: 	lw	%r9, [%r27 + 4]
"00111011011010100000000000000011",	-- 6215: 	lw	%r10, [%r27 + 3]
"00111011011010110000000000000010",	-- 6216: 	lw	%r11, [%r27 + 2]
"00111011011011000000000000000001",	-- 6217: 	lw	%r12, [%r27 + 1]
"00111101001111100000000000000000",	-- 6218: 	sw	%r9, [%sp + 0]
"00111101011111100000000000000001",	-- 6219: 	sw	%r11, [%sp + 1]
"00111101010111100000000000000010",	-- 6220: 	sw	%r10, [%sp + 2]
"00111101100111100000000000000011",	-- 6221: 	sw	%r12, [%sp + 3]
"00111100101111100000000000000100",	-- 6222: 	sw	%r5, [%sp + 4]
"00111100100111100000000000000101",	-- 6223: 	sw	%r4, [%sp + 5]
"00111100111111100000000000000110",	-- 6224: 	sw	%r7, [%sp + 6]
"00111111011111100000000000000111",	-- 6225: 	sw	%r27, [%sp + 7]
"00111101000111100000000000001000",	-- 6226: 	sw	%r8, [%sp + 8]
"00111100011111100000000000001001",	-- 6227: 	sw	%r3, [%sp + 9]
"00111100110111100000000000001010",	-- 6228: 	sw	%r6, [%sp + 10]
"00111100001111100000000000001011",	-- 6229: 	sw	%r1, [%sp + 11]
"00111100010111100000000000001100",	-- 6230: 	sw	%r2, [%sp + 12]
"10000100000000110000100000000000",	-- 6231: 	add	%r1, %r0, %r3
"00111111111111100000000000001101",	-- 6232: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 6233: 	addi	%sp, %sp, 14
"01011000000000000000011010111100",	-- 6234: 	jal	d_vec.2683
"10101011110111100000000000001110",	-- 6235: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 6236: 	lw	%ra, [%sp + 13]
"00111011110000100000000000001011",	-- 6237: 	lw	%r2, [%sp + 11]
"00111011110000110000000000001100",	-- 6238: 	lw	%r3, [%sp + 12]
"10000100011000100010000000000000",	-- 6239: 	add	%r4, %r3, %r2
"00111000100001000000000000000000",	-- 6240: 	lw	%r4, [%r4 + 0]
"11001100000001011111111111111111",	-- 6241: 	lli	%r5, -1
"11001000000001011111111111111111",	-- 6242: 	lhi	%r5, -1
"00101000100001010000000000000010",	-- 6243: 	bneq	%r4, %r5, bneq_else.9124
"01001111111000000000000000000000",	-- 6244: 	jr	%ra
	-- bneq_else.9124:
"00111011110001010000000000001001",	-- 6245: 	lw	%r5, [%sp + 9]
"00111011110110110000000000001010",	-- 6246: 	lw	%r27, [%sp + 10]
"00111100001111100000000000001101",	-- 6247: 	sw	%r1, [%sp + 13]
"00111100100111100000000000001110",	-- 6248: 	sw	%r4, [%sp + 14]
"10000100000001010001000000000000",	-- 6249: 	add	%r2, %r0, %r5
"10000100000001000000100000000000",	-- 6250: 	add	%r1, %r0, %r4
"00111111111111100000000000001111",	-- 6251: 	sw	%ra, [%sp + 15]
"00111011011110100000000000000000",	-- 6252: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010000",	-- 6253: 	addi	%sp, %sp, 16
"01010011010000000000000000000000",	-- 6254: 	jalr	%r26
"10101011110111100000000000010000",	-- 6255: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 6256: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 6257: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 6258: 	bneq	%r1, %r2, bneq_else.9126
"00111011110000010000000000001110",	-- 6259: 	lw	%r1, [%sp + 14]
"00111011110000100000000000001000",	-- 6260: 	lw	%r2, [%sp + 8]
"10000100010000010000100000000000",	-- 6261: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 6262: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001111",	-- 6263: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 6264: 	addi	%sp, %sp, 16
"01011000000000000000011001010110",	-- 6265: 	jal	o_isinvert.2628
"10101011110111100000000000010000",	-- 6266: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 6267: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 6268: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6269: 	bneq	%r1, %r2, bneq_else.9127
"01001111111000000000000000000000",	-- 6270: 	jr	%ra
	-- bneq_else.9127:
"11001100000000010000000000000001",	-- 6271: 	lli	%r1, 1
"00111011110000100000000000001011",	-- 6272: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 6273: 	add	%r1, %r2, %r1
"00111011110000100000000000001100",	-- 6274: 	lw	%r2, [%sp + 12]
"00111011110000110000000000001001",	-- 6275: 	lw	%r3, [%sp + 9]
"00111011110110110000000000000111",	-- 6276: 	lw	%r27, [%sp + 7]
"00111011011110100000000000000000",	-- 6277: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6278: 	jr	%r26
	-- bneq_else.9126:
"11001100000000100000000000000000",	-- 6279: 	lli	%r2, 0
"00111011110000110000000000000110",	-- 6280: 	lw	%r3, [%sp + 6]
"10000100011000100001000000000000",	-- 6281: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 6282: 	lf	%f1, [%r2 + 0]
"00010100000000000000000000000000",	-- 6283: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 6284: 	lhif	%f0, 0.000000
"00111100001111100000000000001111",	-- 6285: 	sw	%r1, [%sp + 15]
"10110000001111100000000000010000",	-- 6286: 	sf	%f1, [%sp + 16]
"00111111111111100000000000010001",	-- 6287: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 6288: 	addi	%sp, %sp, 18
"01011000000000000000010011110011",	-- 6289: 	jal	fless.2532
"10101011110111100000000000010010",	-- 6290: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 6291: 	lw	%ra, [%sp + 17]
"11001100000000100000000000000000",	-- 6292: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6293: 	bneq	%r1, %r2, bneq_else.9129
"01010100000000000001100011101101",	-- 6294: 	j	bneq_cont.9130
	-- bneq_else.9129:
"11001100000000010000000000000000",	-- 6295: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 6296: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 6297: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6298: 	lf	%f1, [%r1 + 0]
"10010011110000000000000000010000",	-- 6299: 	lf	%f0, [%sp + 16]
"00111111111111100000000000010001",	-- 6300: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 6301: 	addi	%sp, %sp, 18
"01011000000000000000010011110011",	-- 6302: 	jal	fless.2532
"10101011110111100000000000010010",	-- 6303: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 6304: 	lw	%ra, [%sp + 17]
"11001100000000100000000000000000",	-- 6305: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6306: 	bneq	%r1, %r2, bneq_else.9131
"01010100000000000001100011101101",	-- 6307: 	j	bneq_cont.9132
	-- bneq_else.9131:
"00010100000000001101011100001010",	-- 6308: 	llif	%f0, 0.010000
"00010000000000000011110000100011",	-- 6309: 	lhif	%f0, 0.010000
"10010011110000010000000000010000",	-- 6310: 	lf	%f1, [%sp + 16]
"11100000001000000000000000000000",	-- 6311: 	addf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 6312: 	lli	%r1, 0
"00111011110000100000000000001101",	-- 6313: 	lw	%r2, [%sp + 13]
"10000100010000010000100000000000",	-- 6314: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6315: 	lf	%f1, [%r1 + 0]
"11101000001000000000100000000000",	-- 6316: 	mulf	%f1, %f1, %f0
"11001100000000010000000000000000",	-- 6317: 	lli	%r1, 0
"00111011110000110000000000000100",	-- 6318: 	lw	%r3, [%sp + 4]
"10000100011000010000100000000000",	-- 6319: 	add	%r1, %r3, %r1
"10010000001000100000000000000000",	-- 6320: 	lf	%f2, [%r1 + 0]
"11100000001000100000100000000000",	-- 6321: 	addf	%f1, %f1, %f2
"11001100000000010000000000000001",	-- 6322: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 6323: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 6324: 	lf	%f2, [%r1 + 0]
"11101000010000000001000000000000",	-- 6325: 	mulf	%f2, %f2, %f0
"11001100000000010000000000000001",	-- 6326: 	lli	%r1, 1
"10000100011000010000100000000000",	-- 6327: 	add	%r1, %r3, %r1
"10010000001000110000000000000000",	-- 6328: 	lf	%f3, [%r1 + 0]
"11100000010000110001000000000000",	-- 6329: 	addf	%f2, %f2, %f3
"11001100000000010000000000000010",	-- 6330: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 6331: 	add	%r1, %r2, %r1
"10010000001000110000000000000000",	-- 6332: 	lf	%f3, [%r1 + 0]
"11101000011000000001100000000000",	-- 6333: 	mulf	%f3, %f3, %f0
"11001100000000010000000000000010",	-- 6334: 	lli	%r1, 2
"10000100011000010000100000000000",	-- 6335: 	add	%r1, %r3, %r1
"10010000001001000000000000000000",	-- 6336: 	lf	%f4, [%r1 + 0]
"11100000011001000001100000000000",	-- 6337: 	addf	%f3, %f3, %f4
"11001100000000010000000000000000",	-- 6338: 	lli	%r1, 0
"00111011110000100000000000001100",	-- 6339: 	lw	%r2, [%sp + 12]
"00111011110110110000000000000011",	-- 6340: 	lw	%r27, [%sp + 3]
"10110000011111100000000000010001",	-- 6341: 	sf	%f3, [%sp + 17]
"10110000010111100000000000010010",	-- 6342: 	sf	%f2, [%sp + 18]
"10110000001111100000000000010011",	-- 6343: 	sf	%f1, [%sp + 19]
"10110000000111100000000000010100",	-- 6344: 	sf	%f0, [%sp + 20]
"00001100001000000000000000000000",	-- 6345: 	movf	%f0, %f1
"00001100010000010000000000000000",	-- 6346: 	movf	%f1, %f2
"00001100011000100000000000000000",	-- 6347: 	movf	%f2, %f3
"00111111111111100000000000010101",	-- 6348: 	sw	%ra, [%sp + 21]
"00111011011110100000000000000000",	-- 6349: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010110",	-- 6350: 	addi	%sp, %sp, 22
"01010011010000000000000000000000",	-- 6351: 	jalr	%r26
"10101011110111100000000000010110",	-- 6352: 	subi	%sp, %sp, 22
"00111011110111110000000000010101",	-- 6353: 	lw	%ra, [%sp + 21]
"11001100000000100000000000000000",	-- 6354: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6355: 	bneq	%r1, %r2, bneq_else.9133
"01010100000000000001100011101101",	-- 6356: 	j	bneq_cont.9134
	-- bneq_else.9133:
"11001100000000010000000000000000",	-- 6357: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 6358: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 6359: 	add	%r1, %r2, %r1
"10010011110000000000000000010100",	-- 6360: 	lf	%f0, [%sp + 20]
"10110000000000010000000000000000",	-- 6361: 	sf	%f0, [%r1 + 0]
"10010011110000000000000000010011",	-- 6362: 	lf	%f0, [%sp + 19]
"10010011110000010000000000010010",	-- 6363: 	lf	%f1, [%sp + 18]
"10010011110000100000000000010001",	-- 6364: 	lf	%f2, [%sp + 17]
"00111011110000010000000000000010",	-- 6365: 	lw	%r1, [%sp + 2]
"00111111111111100000000000010101",	-- 6366: 	sw	%ra, [%sp + 21]
"10100111110111100000000000010110",	-- 6367: 	addi	%sp, %sp, 22
"01011000000000000000010100100110",	-- 6368: 	jal	vecset.2576
"10101011110111100000000000010110",	-- 6369: 	subi	%sp, %sp, 22
"00111011110111110000000000010101",	-- 6370: 	lw	%ra, [%sp + 21]
"11001100000000010000000000000000",	-- 6371: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 6372: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 6373: 	add	%r1, %r2, %r1
"00111011110000100000000000001110",	-- 6374: 	lw	%r2, [%sp + 14]
"00111100010000010000000000000000",	-- 6375: 	sw	%r2, [%r1 + 0]
"11001100000000010000000000000000",	-- 6376: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 6377: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6378: 	add	%r1, %r2, %r1
"00111011110000100000000000001111",	-- 6379: 	lw	%r2, [%sp + 15]
"00111100010000010000000000000000",	-- 6380: 	sw	%r2, [%r1 + 0]
	-- bneq_cont.9134:
	-- bneq_cont.9132:
	-- bneq_cont.9130:
"11001100000000010000000000000001",	-- 6381: 	lli	%r1, 1
"00111011110000100000000000001011",	-- 6382: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 6383: 	add	%r1, %r2, %r1
"00111011110000100000000000001100",	-- 6384: 	lw	%r2, [%sp + 12]
"00111011110000110000000000001001",	-- 6385: 	lw	%r3, [%sp + 9]
"00111011110110110000000000000111",	-- 6386: 	lw	%r27, [%sp + 7]
"00111011011110100000000000000000",	-- 6387: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6388: 	jr	%r26
	-- solve_one_or_network_fast.2872:
"00111011011001000000000000000010",	-- 6389: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 6390: 	lw	%r5, [%r27 + 1]
"10000100010000010011000000000000",	-- 6391: 	add	%r6, %r2, %r1
"00111000110001100000000000000000",	-- 6392: 	lw	%r6, [%r6 + 0]
"11001100000001111111111111111111",	-- 6393: 	lli	%r7, -1
"11001000000001111111111111111111",	-- 6394: 	lhi	%r7, -1
"00101000110001110000000000000010",	-- 6395: 	bneq	%r6, %r7, bneq_else.9135
"01001111111000000000000000000000",	-- 6396: 	jr	%ra
	-- bneq_else.9135:
"10000100101001100010100000000000",	-- 6397: 	add	%r5, %r5, %r6
"00111000101001010000000000000000",	-- 6398: 	lw	%r5, [%r5 + 0]
"11001100000001100000000000000000",	-- 6399: 	lli	%r6, 0
"00111100011111100000000000000000",	-- 6400: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 6401: 	sw	%r2, [%sp + 1]
"00111111011111100000000000000010",	-- 6402: 	sw	%r27, [%sp + 2]
"00111100001111100000000000000011",	-- 6403: 	sw	%r1, [%sp + 3]
"10000100000001010001000000000000",	-- 6404: 	add	%r2, %r0, %r5
"10000100000001100000100000000000",	-- 6405: 	add	%r1, %r0, %r6
"10000100000001001101100000000000",	-- 6406: 	add	%r27, %r0, %r4
"00111111111111100000000000000100",	-- 6407: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 6408: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 6409: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 6410: 	jalr	%r26
"10101011110111100000000000000101",	-- 6411: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6412: 	lw	%ra, [%sp + 4]
"11001100000000010000000000000001",	-- 6413: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 6414: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 6415: 	add	%r1, %r2, %r1
"00111011110000100000000000000001",	-- 6416: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 6417: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000010",	-- 6418: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 6419: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6420: 	jr	%r26
	-- trace_or_matrix_fast.2876:
"00111011011001000000000000000100",	-- 6421: 	lw	%r4, [%r27 + 4]
"00111011011001010000000000000011",	-- 6422: 	lw	%r5, [%r27 + 3]
"00111011011001100000000000000010",	-- 6423: 	lw	%r6, [%r27 + 2]
"00111011011001110000000000000001",	-- 6424: 	lw	%r7, [%r27 + 1]
"10000100010000010100000000000000",	-- 6425: 	add	%r8, %r2, %r1
"00111001000010000000000000000000",	-- 6426: 	lw	%r8, [%r8 + 0]
"11001100000010010000000000000000",	-- 6427: 	lli	%r9, 0
"10000101000010010100100000000000",	-- 6428: 	add	%r9, %r8, %r9
"00111001001010010000000000000000",	-- 6429: 	lw	%r9, [%r9 + 0]
"11001100000010101111111111111111",	-- 6430: 	lli	%r10, -1
"11001000000010101111111111111111",	-- 6431: 	lhi	%r10, -1
"00101001001010100000000000000010",	-- 6432: 	bneq	%r9, %r10, bneq_else.9137
"01001111111000000000000000000000",	-- 6433: 	jr	%ra
	-- bneq_else.9137:
"11001100000010100000000001100011",	-- 6434: 	lli	%r10, 99
"00111100011111100000000000000000",	-- 6435: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 6436: 	sw	%r2, [%sp + 1]
"00111111011111100000000000000010",	-- 6437: 	sw	%r27, [%sp + 2]
"00111100001111100000000000000011",	-- 6438: 	sw	%r1, [%sp + 3]
"00101001001010100000000000001100",	-- 6439: 	bneq	%r9, %r10, bneq_else.9139
"11001100000001000000000000000001",	-- 6440: 	lli	%r4, 1
"10000100000010000001000000000000",	-- 6441: 	add	%r2, %r0, %r8
"10000100000001000000100000000000",	-- 6442: 	add	%r1, %r0, %r4
"10000100000001111101100000000000",	-- 6443: 	add	%r27, %r0, %r7
"00111111111111100000000000000100",	-- 6444: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 6445: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 6446: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 6447: 	jalr	%r26
"10101011110111100000000000000101",	-- 6448: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6449: 	lw	%ra, [%sp + 4]
"01010100000000000001100101011101",	-- 6450: 	j	bneq_cont.9140
	-- bneq_else.9139:
"00111101000111100000000000000100",	-- 6451: 	sw	%r8, [%sp + 4]
"00111100111111100000000000000101",	-- 6452: 	sw	%r7, [%sp + 5]
"00111100100111100000000000000110",	-- 6453: 	sw	%r4, [%sp + 6]
"00111100110111100000000000000111",	-- 6454: 	sw	%r6, [%sp + 7]
"10000100000000110001000000000000",	-- 6455: 	add	%r2, %r0, %r3
"10000100000010010000100000000000",	-- 6456: 	add	%r1, %r0, %r9
"10000100000001011101100000000000",	-- 6457: 	add	%r27, %r0, %r5
"00111111111111100000000000001000",	-- 6458: 	sw	%ra, [%sp + 8]
"00111011011110100000000000000000",	-- 6459: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001001",	-- 6460: 	addi	%sp, %sp, 9
"01010011010000000000000000000000",	-- 6461: 	jalr	%r26
"10101011110111100000000000001001",	-- 6462: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6463: 	lw	%ra, [%sp + 8]
"11001100000000100000000000000000",	-- 6464: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6465: 	bneq	%r1, %r2, bneq_else.9141
"01010100000000000001100101011101",	-- 6466: 	j	bneq_cont.9142
	-- bneq_else.9141:
"11001100000000010000000000000000",	-- 6467: 	lli	%r1, 0
"00111011110000100000000000000111",	-- 6468: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 6469: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 6470: 	lf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 6471: 	lli	%r1, 0
"00111011110000100000000000000110",	-- 6472: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 6473: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6474: 	lf	%f1, [%r1 + 0]
"00111111111111100000000000001000",	-- 6475: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 6476: 	addi	%sp, %sp, 9
"01011000000000000000010011110011",	-- 6477: 	jal	fless.2532
"10101011110111100000000000001001",	-- 6478: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6479: 	lw	%ra, [%sp + 8]
"11001100000000100000000000000000",	-- 6480: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 6481: 	bneq	%r1, %r2, bneq_else.9143
"01010100000000000001100101011101",	-- 6482: 	j	bneq_cont.9144
	-- bneq_else.9143:
"11001100000000010000000000000001",	-- 6483: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 6484: 	lw	%r2, [%sp + 4]
"00111011110000110000000000000000",	-- 6485: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000101",	-- 6486: 	lw	%r27, [%sp + 5]
"00111111111111100000000000001000",	-- 6487: 	sw	%ra, [%sp + 8]
"00111011011110100000000000000000",	-- 6488: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001001",	-- 6489: 	addi	%sp, %sp, 9
"01010011010000000000000000000000",	-- 6490: 	jalr	%r26
"10101011110111100000000000001001",	-- 6491: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6492: 	lw	%ra, [%sp + 8]
	-- bneq_cont.9144:
	-- bneq_cont.9142:
	-- bneq_cont.9140:
"11001100000000010000000000000001",	-- 6493: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 6494: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 6495: 	add	%r1, %r2, %r1
"00111011110000100000000000000001",	-- 6496: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 6497: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000010",	-- 6498: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 6499: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6500: 	jr	%r26
	-- judge_intersection_fast.2880:
"00111011011000100000000000000011",	-- 6501: 	lw	%r2, [%r27 + 3]
"00111011011000110000000000000010",	-- 6502: 	lw	%r3, [%r27 + 2]
"00111011011001000000000000000001",	-- 6503: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 6504: 	lli	%r5, 0
"00010100000000000110101100101000",	-- 6505: 	llif	%f0, 1000000000.000000
"00010000000000000100111001101110",	-- 6506: 	lhif	%f0, 1000000000.000000
"10000100011001010010100000000000",	-- 6507: 	add	%r5, %r3, %r5
"10110000000001010000000000000000",	-- 6508: 	sf	%f0, [%r5 + 0]
"11001100000001010000000000000000",	-- 6509: 	lli	%r5, 0
"11001100000001100000000000000000",	-- 6510: 	lli	%r6, 0
"10000100100001100010000000000000",	-- 6511: 	add	%r4, %r4, %r6
"00111000100001000000000000000000",	-- 6512: 	lw	%r4, [%r4 + 0]
"00111100011111100000000000000000",	-- 6513: 	sw	%r3, [%sp + 0]
"10000100000000010001100000000000",	-- 6514: 	add	%r3, %r0, %r1
"10000100000000101101100000000000",	-- 6515: 	add	%r27, %r0, %r2
"10000100000001000001000000000000",	-- 6516: 	add	%r2, %r0, %r4
"10000100000001010000100000000000",	-- 6517: 	add	%r1, %r0, %r5
"00111111111111100000000000000001",	-- 6518: 	sw	%ra, [%sp + 1]
"00111011011110100000000000000000",	-- 6519: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000010",	-- 6520: 	addi	%sp, %sp, 2
"01010011010000000000000000000000",	-- 6521: 	jalr	%r26
"10101011110111100000000000000010",	-- 6522: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 6523: 	lw	%ra, [%sp + 1]
"11001100000000010000000000000000",	-- 6524: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 6525: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6526: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6527: 	lf	%f1, [%r1 + 0]
"00010100000000001100110011001101",	-- 6528: 	llif	%f0, -0.100000
"00010000000000001011110111001100",	-- 6529: 	lhif	%f0, -0.100000
"10110000001111100000000000000001",	-- 6530: 	sf	%f1, [%sp + 1]
"00111111111111100000000000000010",	-- 6531: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 6532: 	addi	%sp, %sp, 3
"01011000000000000000010011110011",	-- 6533: 	jal	fless.2532
"10101011110111100000000000000011",	-- 6534: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 6535: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000000",	-- 6536: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 6537: 	bneq	%r1, %r2, bneq_else.9145
"11001100000000010000000000000000",	-- 6538: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 6539: 	jr	%ra
	-- bneq_else.9145:
"00010100000000011011110000100000",	-- 6540: 	llif	%f1, 100000000.000000
"00010000000000010100110010111110",	-- 6541: 	lhif	%f1, 100000000.000000
"10010011110000000000000000000001",	-- 6542: 	lf	%f0, [%sp + 1]
"01010100000000000000010011110011",	-- 6543: 	j	fless.2532
	-- get_nvector_rect.2882:
"00111011011000100000000000000010",	-- 6544: 	lw	%r2, [%r27 + 2]
"00111011011000110000000000000001",	-- 6545: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 6546: 	lli	%r4, 0
"10000100011001000001100000000000",	-- 6547: 	add	%r3, %r3, %r4
"00111000011000110000000000000000",	-- 6548: 	lw	%r3, [%r3 + 0]
"00111100010111100000000000000000",	-- 6549: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 6550: 	sw	%r1, [%sp + 1]
"00111100011111100000000000000010",	-- 6551: 	sw	%r3, [%sp + 2]
"10000100000000100000100000000000",	-- 6552: 	add	%r1, %r0, %r2
"00111111111111100000000000000011",	-- 6553: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 6554: 	addi	%sp, %sp, 4
"01011000000000000000010100111010",	-- 6555: 	jal	vecbzero.2584
"10101011110111100000000000000100",	-- 6556: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 6557: 	lw	%ra, [%sp + 3]
"11001100000000010000000000000001",	-- 6558: 	lli	%r1, 1
"00111011110000100000000000000010",	-- 6559: 	lw	%r2, [%sp + 2]
"10001000010000010000100000000000",	-- 6560: 	sub	%r1, %r2, %r1
"11001100000000110000000000000001",	-- 6561: 	lli	%r3, 1
"10001000010000110001000000000000",	-- 6562: 	sub	%r2, %r2, %r3
"00111011110000110000000000000001",	-- 6563: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 6564: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 6565: 	lf	%f0, [%r2 + 0]
"00111100001111100000000000000011",	-- 6566: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 6567: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 6568: 	addi	%sp, %sp, 5
"01011000000000000000010100000010",	-- 6569: 	jal	sgn.2568
"10101011110111100000000000000101",	-- 6570: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6571: 	lw	%ra, [%sp + 4]
"00111111111111100000000000000100",	-- 6572: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 6573: 	addi	%sp, %sp, 5
"01011000000000000010101001010001",	-- 6574: 	jal	yj_fneg
"10101011110111100000000000000101",	-- 6575: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6576: 	lw	%ra, [%sp + 4]
"00111011110000010000000000000011",	-- 6577: 	lw	%r1, [%sp + 3]
"00111011110000100000000000000000",	-- 6578: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6579: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6580: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 6581: 	jr	%ra
	-- get_nvector_plane.2884:
"00111011011000100000000000000001",	-- 6582: 	lw	%r2, [%r27 + 1]
"11001100000000110000000000000000",	-- 6583: 	lli	%r3, 0
"00111100001111100000000000000000",	-- 6584: 	sw	%r1, [%sp + 0]
"00111100011111100000000000000001",	-- 6585: 	sw	%r3, [%sp + 1]
"00111100010111100000000000000010",	-- 6586: 	sw	%r2, [%sp + 2]
"00111111111111100000000000000011",	-- 6587: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 6588: 	addi	%sp, %sp, 4
"01011000000000000000011001011010",	-- 6589: 	jal	o_param_a.2632
"10101011110111100000000000000100",	-- 6590: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 6591: 	lw	%ra, [%sp + 3]
"00111111111111100000000000000011",	-- 6592: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 6593: 	addi	%sp, %sp, 4
"01011000000000000010101001010001",	-- 6594: 	jal	yj_fneg
"10101011110111100000000000000100",	-- 6595: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 6596: 	lw	%ra, [%sp + 3]
"00111011110000010000000000000001",	-- 6597: 	lw	%r1, [%sp + 1]
"00111011110000100000000000000010",	-- 6598: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 6599: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6600: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 6601: 	lli	%r1, 1
"00111011110000110000000000000000",	-- 6602: 	lw	%r3, [%sp + 0]
"00111100001111100000000000000011",	-- 6603: 	sw	%r1, [%sp + 3]
"10000100000000110000100000000000",	-- 6604: 	add	%r1, %r0, %r3
"00111111111111100000000000000100",	-- 6605: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 6606: 	addi	%sp, %sp, 5
"01011000000000000000011001011111",	-- 6607: 	jal	o_param_b.2634
"10101011110111100000000000000101",	-- 6608: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6609: 	lw	%ra, [%sp + 4]
"00111111111111100000000000000100",	-- 6610: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 6611: 	addi	%sp, %sp, 5
"01011000000000000010101001010001",	-- 6612: 	jal	yj_fneg
"10101011110111100000000000000101",	-- 6613: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6614: 	lw	%ra, [%sp + 4]
"00111011110000010000000000000011",	-- 6615: 	lw	%r1, [%sp + 3]
"00111011110000100000000000000010",	-- 6616: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 6617: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6618: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 6619: 	lli	%r1, 2
"00111011110000110000000000000000",	-- 6620: 	lw	%r3, [%sp + 0]
"00111100001111100000000000000100",	-- 6621: 	sw	%r1, [%sp + 4]
"10000100000000110000100000000000",	-- 6622: 	add	%r1, %r0, %r3
"00111111111111100000000000000101",	-- 6623: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 6624: 	addi	%sp, %sp, 6
"01011000000000000000011001100100",	-- 6625: 	jal	o_param_c.2636
"10101011110111100000000000000110",	-- 6626: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 6627: 	lw	%ra, [%sp + 5]
"00111111111111100000000000000101",	-- 6628: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 6629: 	addi	%sp, %sp, 6
"01011000000000000010101001010001",	-- 6630: 	jal	yj_fneg
"10101011110111100000000000000110",	-- 6631: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 6632: 	lw	%ra, [%sp + 5]
"00111011110000010000000000000100",	-- 6633: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000010",	-- 6634: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 6635: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6636: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 6637: 	jr	%ra
	-- get_nvector_second.2886:
"00111011011000100000000000000010",	-- 6638: 	lw	%r2, [%r27 + 2]
"00111011011000110000000000000001",	-- 6639: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 6640: 	lli	%r4, 0
"10000100011001000010000000000000",	-- 6641: 	add	%r4, %r3, %r4
"10010000100000000000000000000000",	-- 6642: 	lf	%f0, [%r4 + 0]
"00111100010111100000000000000000",	-- 6643: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 6644: 	sw	%r1, [%sp + 1]
"00111100011111100000000000000010",	-- 6645: 	sw	%r3, [%sp + 2]
"10110000000111100000000000000011",	-- 6646: 	sf	%f0, [%sp + 3]
"00111111111111100000000000000100",	-- 6647: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 6648: 	addi	%sp, %sp, 5
"01011000000000000000011001101011",	-- 6649: 	jal	o_param_x.2640
"10101011110111100000000000000101",	-- 6650: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 6651: 	lw	%ra, [%sp + 4]
"10010011110000010000000000000011",	-- 6652: 	lf	%f1, [%sp + 3]
"11100100001000000000000000000000",	-- 6653: 	subf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 6654: 	lli	%r1, 1
"00111011110000100000000000000010",	-- 6655: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 6656: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6657: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000001",	-- 6658: 	lw	%r1, [%sp + 1]
"10110000000111100000000000000100",	-- 6659: 	sf	%f0, [%sp + 4]
"10110000001111100000000000000101",	-- 6660: 	sf	%f1, [%sp + 5]
"00111111111111100000000000000110",	-- 6661: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 6662: 	addi	%sp, %sp, 7
"01011000000000000000011001110000",	-- 6663: 	jal	o_param_y.2642
"10101011110111100000000000000111",	-- 6664: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 6665: 	lw	%ra, [%sp + 6]
"10010011110000010000000000000101",	-- 6666: 	lf	%f1, [%sp + 5]
"11100100001000000000000000000000",	-- 6667: 	subf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 6668: 	lli	%r1, 2
"00111011110000100000000000000010",	-- 6669: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 6670: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 6671: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000001",	-- 6672: 	lw	%r1, [%sp + 1]
"10110000000111100000000000000110",	-- 6673: 	sf	%f0, [%sp + 6]
"10110000001111100000000000000111",	-- 6674: 	sf	%f1, [%sp + 7]
"00111111111111100000000000001000",	-- 6675: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 6676: 	addi	%sp, %sp, 9
"01011000000000000000011001110101",	-- 6677: 	jal	o_param_z.2644
"10101011110111100000000000001001",	-- 6678: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6679: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000111",	-- 6680: 	lf	%f1, [%sp + 7]
"11100100001000000000000000000000",	-- 6681: 	subf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6682: 	lw	%r1, [%sp + 1]
"10110000000111100000000000001000",	-- 6683: 	sf	%f0, [%sp + 8]
"00111111111111100000000000001001",	-- 6684: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 6685: 	addi	%sp, %sp, 10
"01011000000000000000011001011010",	-- 6686: 	jal	o_param_a.2632
"10101011110111100000000000001010",	-- 6687: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 6688: 	lw	%ra, [%sp + 9]
"10010011110000010000000000000100",	-- 6689: 	lf	%f1, [%sp + 4]
"11101000001000000000000000000000",	-- 6690: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6691: 	lw	%r1, [%sp + 1]
"10110000000111100000000000001001",	-- 6692: 	sf	%f0, [%sp + 9]
"00111111111111100000000000001010",	-- 6693: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 6694: 	addi	%sp, %sp, 11
"01011000000000000000011001011111",	-- 6695: 	jal	o_param_b.2634
"10101011110111100000000000001011",	-- 6696: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 6697: 	lw	%ra, [%sp + 10]
"10010011110000010000000000000110",	-- 6698: 	lf	%f1, [%sp + 6]
"11101000001000000000000000000000",	-- 6699: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6700: 	lw	%r1, [%sp + 1]
"10110000000111100000000000001010",	-- 6701: 	sf	%f0, [%sp + 10]
"00111111111111100000000000001011",	-- 6702: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 6703: 	addi	%sp, %sp, 12
"01011000000000000000011001100100",	-- 6704: 	jal	o_param_c.2636
"10101011110111100000000000001100",	-- 6705: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 6706: 	lw	%ra, [%sp + 11]
"10010011110000010000000000001000",	-- 6707: 	lf	%f1, [%sp + 8]
"11101000001000000000000000000000",	-- 6708: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6709: 	lw	%r1, [%sp + 1]
"10110000000111100000000000001011",	-- 6710: 	sf	%f0, [%sp + 11]
"00111111111111100000000000001100",	-- 6711: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 6712: 	addi	%sp, %sp, 13
"01011000000000000000011001011000",	-- 6713: 	jal	o_isrot.2630
"10101011110111100000000000001101",	-- 6714: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 6715: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000000",	-- 6716: 	lli	%r2, 0
"00101000001000100000000000001111",	-- 6717: 	bneq	%r1, %r2, bneq_else.9148
"11001100000000010000000000000000",	-- 6718: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 6719: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6720: 	add	%r1, %r2, %r1
"10010011110000000000000000001001",	-- 6721: 	lf	%f0, [%sp + 9]
"10110000000000010000000000000000",	-- 6722: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 6723: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 6724: 	add	%r1, %r2, %r1
"10010011110000000000000000001010",	-- 6725: 	lf	%f0, [%sp + 10]
"10110000000000010000000000000000",	-- 6726: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 6727: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 6728: 	add	%r1, %r2, %r1
"10010011110000000000000000001011",	-- 6729: 	lf	%f0, [%sp + 11]
"10110000000000010000000000000000",	-- 6730: 	sf	%f0, [%r1 + 0]
"01010100000000000001101010101111",	-- 6731: 	j	bneq_cont.9149
	-- bneq_else.9148:
"11001100000000010000000000000000",	-- 6732: 	lli	%r1, 0
"00111011110000100000000000000001",	-- 6733: 	lw	%r2, [%sp + 1]
"00111100001111100000000000001100",	-- 6734: 	sw	%r1, [%sp + 12]
"10000100000000100000100000000000",	-- 6735: 	add	%r1, %r0, %r2
"00111111111111100000000000001101",	-- 6736: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 6737: 	addi	%sp, %sp, 14
"01011000000000000000011010011101",	-- 6738: 	jal	o_param_r3.2660
"10101011110111100000000000001110",	-- 6739: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 6740: 	lw	%ra, [%sp + 13]
"10010011110000010000000000000110",	-- 6741: 	lf	%f1, [%sp + 6]
"11101000001000000000000000000000",	-- 6742: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6743: 	lw	%r1, [%sp + 1]
"10110000000111100000000000001101",	-- 6744: 	sf	%f0, [%sp + 13]
"00111111111111100000000000001110",	-- 6745: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 6746: 	addi	%sp, %sp, 15
"01011000000000000000011010011000",	-- 6747: 	jal	o_param_r2.2658
"10101011110111100000000000001111",	-- 6748: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 6749: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001000",	-- 6750: 	lf	%f1, [%sp + 8]
"11101000001000000000000000000000",	-- 6751: 	mulf	%f0, %f1, %f0
"10010011110000100000000000001101",	-- 6752: 	lf	%f2, [%sp + 13]
"11100000010000000000000000000000",	-- 6753: 	addf	%f0, %f2, %f0
"00111111111111100000000000001110",	-- 6754: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 6755: 	addi	%sp, %sp, 15
"01011000000000000000010011101101",	-- 6756: 	jal	fhalf.2528
"10101011110111100000000000001111",	-- 6757: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 6758: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001001",	-- 6759: 	lf	%f1, [%sp + 9]
"11100000001000000000000000000000",	-- 6760: 	addf	%f0, %f1, %f0
"00111011110000010000000000001100",	-- 6761: 	lw	%r1, [%sp + 12]
"00111011110000100000000000000000",	-- 6762: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6763: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6764: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 6765: 	lli	%r1, 1
"00111011110000110000000000000001",	-- 6766: 	lw	%r3, [%sp + 1]
"00111100001111100000000000001110",	-- 6767: 	sw	%r1, [%sp + 14]
"10000100000000110000100000000000",	-- 6768: 	add	%r1, %r0, %r3
"00111111111111100000000000001111",	-- 6769: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 6770: 	addi	%sp, %sp, 16
"01011000000000000000011010011101",	-- 6771: 	jal	o_param_r3.2660
"10101011110111100000000000010000",	-- 6772: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 6773: 	lw	%ra, [%sp + 15]
"10010011110000010000000000000100",	-- 6774: 	lf	%f1, [%sp + 4]
"11101000001000000000000000000000",	-- 6775: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6776: 	lw	%r1, [%sp + 1]
"10110000000111100000000000001111",	-- 6777: 	sf	%f0, [%sp + 15]
"00111111111111100000000000010000",	-- 6778: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 6779: 	addi	%sp, %sp, 17
"01011000000000000000011010010011",	-- 6780: 	jal	o_param_r1.2656
"10101011110111100000000000010001",	-- 6781: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 6782: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001000",	-- 6783: 	lf	%f1, [%sp + 8]
"11101000001000000000000000000000",	-- 6784: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001111",	-- 6785: 	lf	%f1, [%sp + 15]
"11100000001000000000000000000000",	-- 6786: 	addf	%f0, %f1, %f0
"00111111111111100000000000010000",	-- 6787: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 6788: 	addi	%sp, %sp, 17
"01011000000000000000010011101101",	-- 6789: 	jal	fhalf.2528
"10101011110111100000000000010001",	-- 6790: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 6791: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001010",	-- 6792: 	lf	%f1, [%sp + 10]
"11100000001000000000000000000000",	-- 6793: 	addf	%f0, %f1, %f0
"00111011110000010000000000001110",	-- 6794: 	lw	%r1, [%sp + 14]
"00111011110000100000000000000000",	-- 6795: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6796: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6797: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 6798: 	lli	%r1, 2
"00111011110000110000000000000001",	-- 6799: 	lw	%r3, [%sp + 1]
"00111100001111100000000000010000",	-- 6800: 	sw	%r1, [%sp + 16]
"10000100000000110000100000000000",	-- 6801: 	add	%r1, %r0, %r3
"00111111111111100000000000010001",	-- 6802: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 6803: 	addi	%sp, %sp, 18
"01011000000000000000011010011000",	-- 6804: 	jal	o_param_r2.2658
"10101011110111100000000000010010",	-- 6805: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 6806: 	lw	%ra, [%sp + 17]
"10010011110000010000000000000100",	-- 6807: 	lf	%f1, [%sp + 4]
"11101000001000000000000000000000",	-- 6808: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 6809: 	lw	%r1, [%sp + 1]
"10110000000111100000000000010001",	-- 6810: 	sf	%f0, [%sp + 17]
"00111111111111100000000000010010",	-- 6811: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 6812: 	addi	%sp, %sp, 19
"01011000000000000000011010010011",	-- 6813: 	jal	o_param_r1.2656
"10101011110111100000000000010011",	-- 6814: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 6815: 	lw	%ra, [%sp + 18]
"10010011110000010000000000000110",	-- 6816: 	lf	%f1, [%sp + 6]
"11101000001000000000000000000000",	-- 6817: 	mulf	%f0, %f1, %f0
"10010011110000010000000000010001",	-- 6818: 	lf	%f1, [%sp + 17]
"11100000001000000000000000000000",	-- 6819: 	addf	%f0, %f1, %f0
"00111111111111100000000000010010",	-- 6820: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 6821: 	addi	%sp, %sp, 19
"01011000000000000000010011101101",	-- 6822: 	jal	fhalf.2528
"10101011110111100000000000010011",	-- 6823: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 6824: 	lw	%ra, [%sp + 18]
"10010011110000010000000000001011",	-- 6825: 	lf	%f1, [%sp + 11]
"11100000001000000000000000000000",	-- 6826: 	addf	%f0, %f1, %f0
"00111011110000010000000000010000",	-- 6827: 	lw	%r1, [%sp + 16]
"00111011110000100000000000000000",	-- 6828: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 6829: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6830: 	sf	%f0, [%r1 + 0]
	-- bneq_cont.9149:
"00111011110000010000000000000001",	-- 6831: 	lw	%r1, [%sp + 1]
"00111111111111100000000000010010",	-- 6832: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 6833: 	addi	%sp, %sp, 19
"01011000000000000000011001010110",	-- 6834: 	jal	o_isinvert.2628
"10101011110111100000000000010011",	-- 6835: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 6836: 	lw	%ra, [%sp + 18]
"10000100000000010001000000000000",	-- 6837: 	add	%r2, %r0, %r1
"00111011110000010000000000000000",	-- 6838: 	lw	%r1, [%sp + 0]
"01010100000000000000010101010000",	-- 6839: 	j	vecunit_sgn.2594
	-- get_nvector.2888:
"00111011011000110000000000000011",	-- 6840: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 6841: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 6842: 	lw	%r5, [%r27 + 1]
"00111100011111100000000000000000",	-- 6843: 	sw	%r3, [%sp + 0]
"00111100001111100000000000000001",	-- 6844: 	sw	%r1, [%sp + 1]
"00111100101111100000000000000010",	-- 6845: 	sw	%r5, [%sp + 2]
"00111100010111100000000000000011",	-- 6846: 	sw	%r2, [%sp + 3]
"00111100100111100000000000000100",	-- 6847: 	sw	%r4, [%sp + 4]
"00111111111111100000000000000101",	-- 6848: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 6849: 	addi	%sp, %sp, 6
"01011000000000000000011001010010",	-- 6850: 	jal	o_form.2624
"10101011110111100000000000000110",	-- 6851: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 6852: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000001",	-- 6853: 	lli	%r2, 1
"00101000001000100000000000000101",	-- 6854: 	bneq	%r1, %r2, bneq_else.9150
"00111011110000010000000000000011",	-- 6855: 	lw	%r1, [%sp + 3]
"00111011110110110000000000000100",	-- 6856: 	lw	%r27, [%sp + 4]
"00111011011110100000000000000000",	-- 6857: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6858: 	jr	%r26
	-- bneq_else.9150:
"11001100000000100000000000000010",	-- 6859: 	lli	%r2, 2
"00101000001000100000000000000101",	-- 6860: 	bneq	%r1, %r2, bneq_else.9151
"00111011110000010000000000000001",	-- 6861: 	lw	%r1, [%sp + 1]
"00111011110110110000000000000010",	-- 6862: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 6863: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6864: 	jr	%r26
	-- bneq_else.9151:
"00111011110000010000000000000001",	-- 6865: 	lw	%r1, [%sp + 1]
"00111011110110110000000000000000",	-- 6866: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 6867: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 6868: 	jr	%r26
	-- utexture.2891:
"00111011011000110000000000000001",	-- 6869: 	lw	%r3, [%r27 + 1]
"00111100010111100000000000000000",	-- 6870: 	sw	%r2, [%sp + 0]
"00111100011111100000000000000001",	-- 6871: 	sw	%r3, [%sp + 1]
"00111100001111100000000000000010",	-- 6872: 	sw	%r1, [%sp + 2]
"00111111111111100000000000000011",	-- 6873: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 6874: 	addi	%sp, %sp, 4
"01011000000000000000011001010000",	-- 6875: 	jal	o_texturetype.2622
"10101011110111100000000000000100",	-- 6876: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 6877: 	lw	%ra, [%sp + 3]
"11001100000000100000000000000000",	-- 6878: 	lli	%r2, 0
"00111011110000110000000000000010",	-- 6879: 	lw	%r3, [%sp + 2]
"00111100001111100000000000000011",	-- 6880: 	sw	%r1, [%sp + 3]
"00111100010111100000000000000100",	-- 6881: 	sw	%r2, [%sp + 4]
"10000100000000110000100000000000",	-- 6882: 	add	%r1, %r0, %r3
"00111111111111100000000000000101",	-- 6883: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 6884: 	addi	%sp, %sp, 6
"01011000000000000000011010000100",	-- 6885: 	jal	o_color_red.2650
"10101011110111100000000000000110",	-- 6886: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 6887: 	lw	%ra, [%sp + 5]
"00111011110000010000000000000100",	-- 6888: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000001",	-- 6889: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 6890: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6891: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 6892: 	lli	%r1, 1
"00111011110000110000000000000010",	-- 6893: 	lw	%r3, [%sp + 2]
"00111100001111100000000000000101",	-- 6894: 	sw	%r1, [%sp + 5]
"10000100000000110000100000000000",	-- 6895: 	add	%r1, %r0, %r3
"00111111111111100000000000000110",	-- 6896: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 6897: 	addi	%sp, %sp, 7
"01011000000000000000011010001001",	-- 6898: 	jal	o_color_green.2652
"10101011110111100000000000000111",	-- 6899: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 6900: 	lw	%ra, [%sp + 6]
"00111011110000010000000000000101",	-- 6901: 	lw	%r1, [%sp + 5]
"00111011110000100000000000000001",	-- 6902: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 6903: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6904: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000010",	-- 6905: 	lli	%r1, 2
"00111011110000110000000000000010",	-- 6906: 	lw	%r3, [%sp + 2]
"00111100001111100000000000000110",	-- 6907: 	sw	%r1, [%sp + 6]
"10000100000000110000100000000000",	-- 6908: 	add	%r1, %r0, %r3
"00111111111111100000000000000111",	-- 6909: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 6910: 	addi	%sp, %sp, 8
"01011000000000000000011010001110",	-- 6911: 	jal	o_color_blue.2654
"10101011110111100000000000001000",	-- 6912: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 6913: 	lw	%ra, [%sp + 7]
"00111011110000010000000000000110",	-- 6914: 	lw	%r1, [%sp + 6]
"00111011110000100000000000000001",	-- 6915: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 6916: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 6917: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000001",	-- 6918: 	lli	%r1, 1
"00111011110000110000000000000011",	-- 6919: 	lw	%r3, [%sp + 3]
"00101000011000010000000001100000",	-- 6920: 	bneq	%r3, %r1, bneq_else.9152
"11001100000000010000000000000000",	-- 6921: 	lli	%r1, 0
"00111011110000110000000000000000",	-- 6922: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 6923: 	add	%r1, %r3, %r1
"10010000001000000000000000000000",	-- 6924: 	lf	%f0, [%r1 + 0]
"00111011110000010000000000000010",	-- 6925: 	lw	%r1, [%sp + 2]
"10110000000111100000000000000111",	-- 6926: 	sf	%f0, [%sp + 7]
"00111111111111100000000000001000",	-- 6927: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 6928: 	addi	%sp, %sp, 9
"01011000000000000000011001101011",	-- 6929: 	jal	o_param_x.2640
"10101011110111100000000000001001",	-- 6930: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 6931: 	lw	%ra, [%sp + 8]
"10010011110000010000000000000111",	-- 6932: 	lf	%f1, [%sp + 7]
"11100100001000000000000000000000",	-- 6933: 	subf	%f0, %f1, %f0
"00010100000000011100110011001101",	-- 6934: 	llif	%f1, 0.050000
"00010000000000010011110101001100",	-- 6935: 	lhif	%f1, 0.050000
"11101000000000010000100000000000",	-- 6936: 	mulf	%f1, %f0, %f1
"10110000000111100000000000001000",	-- 6937: 	sf	%f0, [%sp + 8]
"00001100001000000000000000000000",	-- 6938: 	movf	%f0, %f1
"00111111111111100000000000001001",	-- 6939: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 6940: 	addi	%sp, %sp, 10
"01011000000000000010101000110010",	-- 6941: 	jal	yj_floor
"10101011110111100000000000001010",	-- 6942: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 6943: 	lw	%ra, [%sp + 9]
"00010100000000010000000000000000",	-- 6944: 	llif	%f1, 20.000000
"00010000000000010100000110100000",	-- 6945: 	lhif	%f1, 20.000000
"11101000000000010000000000000000",	-- 6946: 	mulf	%f0, %f0, %f1
"10010011110000010000000000001000",	-- 6947: 	lf	%f1, [%sp + 8]
"11100100001000000000000000000000",	-- 6948: 	subf	%f0, %f1, %f0
"00010100000000010000000000000000",	-- 6949: 	llif	%f1, 10.000000
"00010000000000010100000100100000",	-- 6950: 	lhif	%f1, 10.000000
"00111111111111100000000000001001",	-- 6951: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 6952: 	addi	%sp, %sp, 10
"01011000000000000000010011110011",	-- 6953: 	jal	fless.2532
"10101011110111100000000000001010",	-- 6954: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 6955: 	lw	%ra, [%sp + 9]
"11001100000000100000000000000010",	-- 6956: 	lli	%r2, 2
"00111011110000110000000000000000",	-- 6957: 	lw	%r3, [%sp + 0]
"10000100011000100001000000000000",	-- 6958: 	add	%r2, %r3, %r2
"10010000010000000000000000000000",	-- 6959: 	lf	%f0, [%r2 + 0]
"00111011110000100000000000000010",	-- 6960: 	lw	%r2, [%sp + 2]
"00111100001111100000000000001001",	-- 6961: 	sw	%r1, [%sp + 9]
"10110000000111100000000000001010",	-- 6962: 	sf	%f0, [%sp + 10]
"10000100000000100000100000000000",	-- 6963: 	add	%r1, %r0, %r2
"00111111111111100000000000001011",	-- 6964: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 6965: 	addi	%sp, %sp, 12
"01011000000000000000011001110101",	-- 6966: 	jal	o_param_z.2644
"10101011110111100000000000001100",	-- 6967: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 6968: 	lw	%ra, [%sp + 11]
"10010011110000010000000000001010",	-- 6969: 	lf	%f1, [%sp + 10]
"11100100001000000000000000000000",	-- 6970: 	subf	%f0, %f1, %f0
"00010100000000011100110011001101",	-- 6971: 	llif	%f1, 0.050000
"00010000000000010011110101001100",	-- 6972: 	lhif	%f1, 0.050000
"11101000000000010000100000000000",	-- 6973: 	mulf	%f1, %f0, %f1
"10110000000111100000000000001011",	-- 6974: 	sf	%f0, [%sp + 11]
"00001100001000000000000000000000",	-- 6975: 	movf	%f0, %f1
"00111111111111100000000000001100",	-- 6976: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 6977: 	addi	%sp, %sp, 13
"01011000000000000010101000110010",	-- 6978: 	jal	yj_floor
"10101011110111100000000000001101",	-- 6979: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 6980: 	lw	%ra, [%sp + 12]
"00010100000000010000000000000000",	-- 6981: 	llif	%f1, 20.000000
"00010000000000010100000110100000",	-- 6982: 	lhif	%f1, 20.000000
"11101000000000010000000000000000",	-- 6983: 	mulf	%f0, %f0, %f1
"10010011110000010000000000001011",	-- 6984: 	lf	%f1, [%sp + 11]
"11100100001000000000000000000000",	-- 6985: 	subf	%f0, %f1, %f0
"00010100000000010000000000000000",	-- 6986: 	llif	%f1, 10.000000
"00010000000000010100000100100000",	-- 6987: 	lhif	%f1, 10.000000
"00111111111111100000000000001100",	-- 6988: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 6989: 	addi	%sp, %sp, 13
"01011000000000000000010011110011",	-- 6990: 	jal	fless.2532
"10101011110111100000000000001101",	-- 6991: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 6992: 	lw	%ra, [%sp + 12]
"11001100000000100000000000000001",	-- 6993: 	lli	%r2, 1
"11001100000000110000000000000000",	-- 6994: 	lli	%r3, 0
"00111011110001000000000000001001",	-- 6995: 	lw	%r4, [%sp + 9]
"00101000100000110000000000001001",	-- 6996: 	bneq	%r4, %r3, bneq_else.9153
"11001100000000110000000000000000",	-- 6997: 	lli	%r3, 0
"00101000001000110000000000000100",	-- 6998: 	bneq	%r1, %r3, bneq_else.9155
"00010100000000000000000000000000",	-- 6999: 	llif	%f0, 255.000000
"00010000000000000100001101111111",	-- 7000: 	lhif	%f0, 255.000000
"01010100000000000001101101011100",	-- 7001: 	j	bneq_cont.9156
	-- bneq_else.9155:
"00010100000000000000000000000000",	-- 7002: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 7003: 	lhif	%f0, 0.000000
	-- bneq_cont.9156:
"01010100000000000001101101100100",	-- 7004: 	j	bneq_cont.9154
	-- bneq_else.9153:
"11001100000000110000000000000000",	-- 7005: 	lli	%r3, 0
"00101000001000110000000000000100",	-- 7006: 	bneq	%r1, %r3, bneq_else.9157
"00010100000000000000000000000000",	-- 7007: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 7008: 	lhif	%f0, 0.000000
"01010100000000000001101101100100",	-- 7009: 	j	bneq_cont.9158
	-- bneq_else.9157:
"00010100000000000000000000000000",	-- 7010: 	llif	%f0, 255.000000
"00010000000000000100001101111111",	-- 7011: 	lhif	%f0, 255.000000
	-- bneq_cont.9158:
	-- bneq_cont.9154:
"00111011110000010000000000000001",	-- 7012: 	lw	%r1, [%sp + 1]
"10000100001000100000100000000000",	-- 7013: 	add	%r1, %r1, %r2
"10110000000000010000000000000000",	-- 7014: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 7015: 	jr	%ra
	-- bneq_else.9152:
"11001100000000010000000000000010",	-- 7016: 	lli	%r1, 2
"00101000011000010000000000100011",	-- 7017: 	bneq	%r3, %r1, bneq_else.9160
"11001100000000010000000000000001",	-- 7018: 	lli	%r1, 1
"00111011110000110000000000000000",	-- 7019: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 7020: 	add	%r1, %r3, %r1
"10010000001000000000000000000000",	-- 7021: 	lf	%f0, [%r1 + 0]
"00010100000000010000000000000000",	-- 7022: 	llif	%f1, 0.250000
"00010000000000010011111010000000",	-- 7023: 	lhif	%f1, 0.250000
"11101000000000010000000000000000",	-- 7024: 	mulf	%f0, %f0, %f1
"00111111111111100000000000001100",	-- 7025: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 7026: 	addi	%sp, %sp, 13
"01011000000000000000010001011001",	-- 7027: 	jal	sin.2516
"10101011110111100000000000001101",	-- 7028: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 7029: 	lw	%ra, [%sp + 12]
"00111111111111100000000000001100",	-- 7030: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 7031: 	addi	%sp, %sp, 13
"01011000000000000000010011110001",	-- 7032: 	jal	fsqr.2530
"10101011110111100000000000001101",	-- 7033: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 7034: 	lw	%ra, [%sp + 12]
"11001100000000010000000000000000",	-- 7035: 	lli	%r1, 0
"00010100000000010000000000000000",	-- 7036: 	llif	%f1, 255.000000
"00010000000000010100001101111111",	-- 7037: 	lhif	%f1, 255.000000
"11101000001000000000100000000000",	-- 7038: 	mulf	%f1, %f1, %f0
"00111011110000100000000000000001",	-- 7039: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 7040: 	add	%r1, %r2, %r1
"10110000001000010000000000000000",	-- 7041: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000001",	-- 7042: 	lli	%r1, 1
"00010100000000010000000000000000",	-- 7043: 	llif	%f1, 255.000000
"00010000000000010100001101111111",	-- 7044: 	lhif	%f1, 255.000000
"00010100000000100000000000000000",	-- 7045: 	llif	%f2, 1.000000
"00010000000000100011111110000000",	-- 7046: 	lhif	%f2, 1.000000
"11100100010000000000000000000000",	-- 7047: 	subf	%f0, %f2, %f0
"11101000001000000000000000000000",	-- 7048: 	mulf	%f0, %f1, %f0
"10000100010000010000100000000000",	-- 7049: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 7050: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 7051: 	jr	%ra
	-- bneq_else.9160:
"11001100000000010000000000000011",	-- 7052: 	lli	%r1, 3
"00101000011000010000000001011100",	-- 7053: 	bneq	%r3, %r1, bneq_else.9162
"11001100000000010000000000000000",	-- 7054: 	lli	%r1, 0
"00111011110000110000000000000000",	-- 7055: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 7056: 	add	%r1, %r3, %r1
"10010000001000000000000000000000",	-- 7057: 	lf	%f0, [%r1 + 0]
"00111011110000010000000000000010",	-- 7058: 	lw	%r1, [%sp + 2]
"10110000000111100000000000001100",	-- 7059: 	sf	%f0, [%sp + 12]
"00111111111111100000000000001101",	-- 7060: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 7061: 	addi	%sp, %sp, 14
"01011000000000000000011001101011",	-- 7062: 	jal	o_param_x.2640
"10101011110111100000000000001110",	-- 7063: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 7064: 	lw	%ra, [%sp + 13]
"10010011110000010000000000001100",	-- 7065: 	lf	%f1, [%sp + 12]
"11100100001000000000000000000000",	-- 7066: 	subf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 7067: 	lli	%r1, 2
"00111011110000100000000000000000",	-- 7068: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 7069: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 7070: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000010",	-- 7071: 	lw	%r1, [%sp + 2]
"10110000000111100000000000001101",	-- 7072: 	sf	%f0, [%sp + 13]
"10110000001111100000000000001110",	-- 7073: 	sf	%f1, [%sp + 14]
"00111111111111100000000000001111",	-- 7074: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 7075: 	addi	%sp, %sp, 16
"01011000000000000000011001110101",	-- 7076: 	jal	o_param_z.2644
"10101011110111100000000000010000",	-- 7077: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 7078: 	lw	%ra, [%sp + 15]
"10010011110000010000000000001110",	-- 7079: 	lf	%f1, [%sp + 14]
"11100100001000000000000000000000",	-- 7080: 	subf	%f0, %f1, %f0
"10010011110000010000000000001101",	-- 7081: 	lf	%f1, [%sp + 13]
"10110000000111100000000000001111",	-- 7082: 	sf	%f0, [%sp + 15]
"00001100001000000000000000000000",	-- 7083: 	movf	%f0, %f1
"00111111111111100000000000010000",	-- 7084: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 7085: 	addi	%sp, %sp, 17
"01011000000000000000010011110001",	-- 7086: 	jal	fsqr.2530
"10101011110111100000000000010001",	-- 7087: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 7088: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001111",	-- 7089: 	lf	%f1, [%sp + 15]
"10110000000111100000000000010000",	-- 7090: 	sf	%f0, [%sp + 16]
"00001100001000000000000000000000",	-- 7091: 	movf	%f0, %f1
"00111111111111100000000000010001",	-- 7092: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 7093: 	addi	%sp, %sp, 18
"01011000000000000000010011110001",	-- 7094: 	jal	fsqr.2530
"10101011110111100000000000010010",	-- 7095: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 7096: 	lw	%ra, [%sp + 17]
"10010011110000010000000000010000",	-- 7097: 	lf	%f1, [%sp + 16]
"11100000001000000000000000000000",	-- 7098: 	addf	%f0, %f1, %f0
"00111111111111100000000000010001",	-- 7099: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 7100: 	addi	%sp, %sp, 18
"01011000000000000010101000110000",	-- 7101: 	jal	yj_sqrt
"10101011110111100000000000010010",	-- 7102: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 7103: 	lw	%ra, [%sp + 17]
"00010100000000010000000000000000",	-- 7104: 	llif	%f1, 10.000000
"00010000000000010100000100100000",	-- 7105: 	lhif	%f1, 10.000000
"11101100000000010000000000000000",	-- 7106: 	divf	%f0, %f0, %f1
"10110000000111100000000000010001",	-- 7107: 	sf	%f0, [%sp + 17]
"00111111111111100000000000010010",	-- 7108: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 7109: 	addi	%sp, %sp, 19
"01011000000000000010101000110010",	-- 7110: 	jal	yj_floor
"10101011110111100000000000010011",	-- 7111: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 7112: 	lw	%ra, [%sp + 18]
"10010011110000010000000000010001",	-- 7113: 	lf	%f1, [%sp + 17]
"11100100001000000000000000000000",	-- 7114: 	subf	%f0, %f1, %f0
"00010100000000010000111111011100",	-- 7115: 	llif	%f1, 3.141593
"00010000000000010100000001001001",	-- 7116: 	lhif	%f1, 3.141593
"11101000000000010000000000000000",	-- 7117: 	mulf	%f0, %f0, %f1
"00111111111111100000000000010010",	-- 7118: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 7119: 	addi	%sp, %sp, 19
"01011000000000000000010010011000",	-- 7120: 	jal	cos.2518
"10101011110111100000000000010011",	-- 7121: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 7122: 	lw	%ra, [%sp + 18]
"00111111111111100000000000010010",	-- 7123: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 7124: 	addi	%sp, %sp, 19
"01011000000000000000010011110001",	-- 7125: 	jal	fsqr.2530
"10101011110111100000000000010011",	-- 7126: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 7127: 	lw	%ra, [%sp + 18]
"11001100000000010000000000000001",	-- 7128: 	lli	%r1, 1
"00010100000000010000000000000000",	-- 7129: 	llif	%f1, 255.000000
"00010000000000010100001101111111",	-- 7130: 	lhif	%f1, 255.000000
"11101000000000010000100000000000",	-- 7131: 	mulf	%f1, %f0, %f1
"00111011110000100000000000000001",	-- 7132: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 7133: 	add	%r1, %r2, %r1
"10110000001000010000000000000000",	-- 7134: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 7135: 	lli	%r1, 2
"00010100000000010000000000000000",	-- 7136: 	llif	%f1, 1.000000
"00010000000000010011111110000000",	-- 7137: 	lhif	%f1, 1.000000
"11100100001000000000000000000000",	-- 7138: 	subf	%f0, %f1, %f0
"00010100000000010000000000000000",	-- 7139: 	llif	%f1, 255.000000
"00010000000000010100001101111111",	-- 7140: 	lhif	%f1, 255.000000
"11101000000000010000000000000000",	-- 7141: 	mulf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 7142: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 7143: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 7144: 	jr	%ra
	-- bneq_else.9162:
"11001100000000010000000000000100",	-- 7145: 	lli	%r1, 4
"00101000011000010000000011111000",	-- 7146: 	bneq	%r3, %r1, bneq_else.9164
"11001100000000010000000000000000",	-- 7147: 	lli	%r1, 0
"00111011110000110000000000000000",	-- 7148: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 7149: 	add	%r1, %r3, %r1
"10010000001000000000000000000000",	-- 7150: 	lf	%f0, [%r1 + 0]
"00111011110000010000000000000010",	-- 7151: 	lw	%r1, [%sp + 2]
"10110000000111100000000000010010",	-- 7152: 	sf	%f0, [%sp + 18]
"00111111111111100000000000010011",	-- 7153: 	sw	%ra, [%sp + 19]
"10100111110111100000000000010100",	-- 7154: 	addi	%sp, %sp, 20
"01011000000000000000011001101011",	-- 7155: 	jal	o_param_x.2640
"10101011110111100000000000010100",	-- 7156: 	subi	%sp, %sp, 20
"00111011110111110000000000010011",	-- 7157: 	lw	%ra, [%sp + 19]
"10010011110000010000000000010010",	-- 7158: 	lf	%f1, [%sp + 18]
"11100100001000000000000000000000",	-- 7159: 	subf	%f0, %f1, %f0
"00111011110000010000000000000010",	-- 7160: 	lw	%r1, [%sp + 2]
"10110000000111100000000000010011",	-- 7161: 	sf	%f0, [%sp + 19]
"00111111111111100000000000010100",	-- 7162: 	sw	%ra, [%sp + 20]
"10100111110111100000000000010101",	-- 7163: 	addi	%sp, %sp, 21
"01011000000000000000011001011010",	-- 7164: 	jal	o_param_a.2632
"10101011110111100000000000010101",	-- 7165: 	subi	%sp, %sp, 21
"00111011110111110000000000010100",	-- 7166: 	lw	%ra, [%sp + 20]
"00111111111111100000000000010100",	-- 7167: 	sw	%ra, [%sp + 20]
"10100111110111100000000000010101",	-- 7168: 	addi	%sp, %sp, 21
"01011000000000000010101000110000",	-- 7169: 	jal	yj_sqrt
"10101011110111100000000000010101",	-- 7170: 	subi	%sp, %sp, 21
"00111011110111110000000000010100",	-- 7171: 	lw	%ra, [%sp + 20]
"10010011110000010000000000010011",	-- 7172: 	lf	%f1, [%sp + 19]
"11101000001000000000000000000000",	-- 7173: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000010",	-- 7174: 	lli	%r1, 2
"00111011110000100000000000000000",	-- 7175: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 7176: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 7177: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000010",	-- 7178: 	lw	%r1, [%sp + 2]
"10110000000111100000000000010100",	-- 7179: 	sf	%f0, [%sp + 20]
"10110000001111100000000000010101",	-- 7180: 	sf	%f1, [%sp + 21]
"00111111111111100000000000010110",	-- 7181: 	sw	%ra, [%sp + 22]
"10100111110111100000000000010111",	-- 7182: 	addi	%sp, %sp, 23
"01011000000000000000011001110101",	-- 7183: 	jal	o_param_z.2644
"10101011110111100000000000010111",	-- 7184: 	subi	%sp, %sp, 23
"00111011110111110000000000010110",	-- 7185: 	lw	%ra, [%sp + 22]
"10010011110000010000000000010101",	-- 7186: 	lf	%f1, [%sp + 21]
"11100100001000000000000000000000",	-- 7187: 	subf	%f0, %f1, %f0
"00111011110000010000000000000010",	-- 7188: 	lw	%r1, [%sp + 2]
"10110000000111100000000000010110",	-- 7189: 	sf	%f0, [%sp + 22]
"00111111111111100000000000010111",	-- 7190: 	sw	%ra, [%sp + 23]
"10100111110111100000000000011000",	-- 7191: 	addi	%sp, %sp, 24
"01011000000000000000011001100100",	-- 7192: 	jal	o_param_c.2636
"10101011110111100000000000011000",	-- 7193: 	subi	%sp, %sp, 24
"00111011110111110000000000010111",	-- 7194: 	lw	%ra, [%sp + 23]
"00111111111111100000000000010111",	-- 7195: 	sw	%ra, [%sp + 23]
"10100111110111100000000000011000",	-- 7196: 	addi	%sp, %sp, 24
"01011000000000000010101000110000",	-- 7197: 	jal	yj_sqrt
"10101011110111100000000000011000",	-- 7198: 	subi	%sp, %sp, 24
"00111011110111110000000000010111",	-- 7199: 	lw	%ra, [%sp + 23]
"10010011110000010000000000010110",	-- 7200: 	lf	%f1, [%sp + 22]
"11101000001000000000000000000000",	-- 7201: 	mulf	%f0, %f1, %f0
"10010011110000010000000000010100",	-- 7202: 	lf	%f1, [%sp + 20]
"10110000000111100000000000010111",	-- 7203: 	sf	%f0, [%sp + 23]
"00001100001000000000000000000000",	-- 7204: 	movf	%f0, %f1
"00111111111111100000000000011000",	-- 7205: 	sw	%ra, [%sp + 24]
"10100111110111100000000000011001",	-- 7206: 	addi	%sp, %sp, 25
"01011000000000000000010011110001",	-- 7207: 	jal	fsqr.2530
"10101011110111100000000000011001",	-- 7208: 	subi	%sp, %sp, 25
"00111011110111110000000000011000",	-- 7209: 	lw	%ra, [%sp + 24]
"10010011110000010000000000010111",	-- 7210: 	lf	%f1, [%sp + 23]
"10110000000111100000000000011000",	-- 7211: 	sf	%f0, [%sp + 24]
"00001100001000000000000000000000",	-- 7212: 	movf	%f0, %f1
"00111111111111100000000000011001",	-- 7213: 	sw	%ra, [%sp + 25]
"10100111110111100000000000011010",	-- 7214: 	addi	%sp, %sp, 26
"01011000000000000000010011110001",	-- 7215: 	jal	fsqr.2530
"10101011110111100000000000011010",	-- 7216: 	subi	%sp, %sp, 26
"00111011110111110000000000011001",	-- 7217: 	lw	%ra, [%sp + 25]
"10010011110000010000000000011000",	-- 7218: 	lf	%f1, [%sp + 24]
"11100000001000000000000000000000",	-- 7219: 	addf	%f0, %f1, %f0
"10010011110000010000000000010100",	-- 7220: 	lf	%f1, [%sp + 20]
"10110000000111100000000000011001",	-- 7221: 	sf	%f0, [%sp + 25]
"00001100001000000000000000000000",	-- 7222: 	movf	%f0, %f1
"00111111111111100000000000011010",	-- 7223: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 7224: 	addi	%sp, %sp, 27
"01011000000000000010101001001111",	-- 7225: 	jal	yj_fabs
"10101011110111100000000000011011",	-- 7226: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 7227: 	lw	%ra, [%sp + 26]
"00010100000000011011011100010111",	-- 7228: 	llif	%f1, 0.000100
"00010000000000010011100011010001",	-- 7229: 	lhif	%f1, 0.000100
"00111111111111100000000000011010",	-- 7230: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 7231: 	addi	%sp, %sp, 27
"01011000000000000000010011110011",	-- 7232: 	jal	fless.2532
"10101011110111100000000000011011",	-- 7233: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 7234: 	lw	%ra, [%sp + 26]
"11001100000000100000000000000000",	-- 7235: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 7236: 	bneq	%r1, %r2, bneq_else.9165
"10010011110000000000000000010100",	-- 7237: 	lf	%f0, [%sp + 20]
"10010011110000010000000000010111",	-- 7238: 	lf	%f1, [%sp + 23]
"11101100001000000000000000000000",	-- 7239: 	divf	%f0, %f1, %f0
"00111111111111100000000000011010",	-- 7240: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 7241: 	addi	%sp, %sp, 27
"01011000000000000010101001001111",	-- 7242: 	jal	yj_fabs
"10101011110111100000000000011011",	-- 7243: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 7244: 	lw	%ra, [%sp + 26]
"00111111111111100000000000011010",	-- 7245: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 7246: 	addi	%sp, %sp, 27
"01011000000000000000010010011110",	-- 7247: 	jal	atan.2520
"10101011110111100000000000011011",	-- 7248: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 7249: 	lw	%ra, [%sp + 26]
"00010100000000010000000000000000",	-- 7250: 	llif	%f1, 30.000000
"00010000000000010100000111110000",	-- 7251: 	lhif	%f1, 30.000000
"11101000000000010000000000000000",	-- 7252: 	mulf	%f0, %f0, %f1
"00010100000000010000111111011100",	-- 7253: 	llif	%f1, 3.141593
"00010000000000010100000001001001",	-- 7254: 	lhif	%f1, 3.141593
"11101100000000010000000000000000",	-- 7255: 	divf	%f0, %f0, %f1
"01010100000000000001110001011011",	-- 7256: 	j	bneq_cont.9166
	-- bneq_else.9165:
"00010100000000000000000000000000",	-- 7257: 	llif	%f0, 15.000000
"00010000000000000100000101110000",	-- 7258: 	lhif	%f0, 15.000000
	-- bneq_cont.9166:
"10110000000111100000000000011010",	-- 7259: 	sf	%f0, [%sp + 26]
"00111111111111100000000000011011",	-- 7260: 	sw	%ra, [%sp + 27]
"10100111110111100000000000011100",	-- 7261: 	addi	%sp, %sp, 28
"01011000000000000010101000110010",	-- 7262: 	jal	yj_floor
"10101011110111100000000000011100",	-- 7263: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 7264: 	lw	%ra, [%sp + 27]
"10010011110000010000000000011010",	-- 7265: 	lf	%f1, [%sp + 26]
"11100100001000000000000000000000",	-- 7266: 	subf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 7267: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 7268: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 7269: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 7270: 	lf	%f1, [%r1 + 0]
"00111011110000010000000000000010",	-- 7271: 	lw	%r1, [%sp + 2]
"10110000000111100000000000011011",	-- 7272: 	sf	%f0, [%sp + 27]
"10110000001111100000000000011100",	-- 7273: 	sf	%f1, [%sp + 28]
"00111111111111100000000000011101",	-- 7274: 	sw	%ra, [%sp + 29]
"10100111110111100000000000011110",	-- 7275: 	addi	%sp, %sp, 30
"01011000000000000000011001110000",	-- 7276: 	jal	o_param_y.2642
"10101011110111100000000000011110",	-- 7277: 	subi	%sp, %sp, 30
"00111011110111110000000000011101",	-- 7278: 	lw	%ra, [%sp + 29]
"10010011110000010000000000011100",	-- 7279: 	lf	%f1, [%sp + 28]
"11100100001000000000000000000000",	-- 7280: 	subf	%f0, %f1, %f0
"00111011110000010000000000000010",	-- 7281: 	lw	%r1, [%sp + 2]
"10110000000111100000000000011101",	-- 7282: 	sf	%f0, [%sp + 29]
"00111111111111100000000000011110",	-- 7283: 	sw	%ra, [%sp + 30]
"10100111110111100000000000011111",	-- 7284: 	addi	%sp, %sp, 31
"01011000000000000000011001011111",	-- 7285: 	jal	o_param_b.2634
"10101011110111100000000000011111",	-- 7286: 	subi	%sp, %sp, 31
"00111011110111110000000000011110",	-- 7287: 	lw	%ra, [%sp + 30]
"00111111111111100000000000011110",	-- 7288: 	sw	%ra, [%sp + 30]
"10100111110111100000000000011111",	-- 7289: 	addi	%sp, %sp, 31
"01011000000000000010101000110000",	-- 7290: 	jal	yj_sqrt
"10101011110111100000000000011111",	-- 7291: 	subi	%sp, %sp, 31
"00111011110111110000000000011110",	-- 7292: 	lw	%ra, [%sp + 30]
"10010011110000010000000000011101",	-- 7293: 	lf	%f1, [%sp + 29]
"11101000001000000000000000000000",	-- 7294: 	mulf	%f0, %f1, %f0
"10010011110000010000000000011001",	-- 7295: 	lf	%f1, [%sp + 25]
"10110000000111100000000000011110",	-- 7296: 	sf	%f0, [%sp + 30]
"00001100001000000000000000000000",	-- 7297: 	movf	%f0, %f1
"00111111111111100000000000011111",	-- 7298: 	sw	%ra, [%sp + 31]
"10100111110111100000000000100000",	-- 7299: 	addi	%sp, %sp, 32
"01011000000000000010101001001111",	-- 7300: 	jal	yj_fabs
"10101011110111100000000000100000",	-- 7301: 	subi	%sp, %sp, 32
"00111011110111110000000000011111",	-- 7302: 	lw	%ra, [%sp + 31]
"00010100000000011011011100010111",	-- 7303: 	llif	%f1, 0.000100
"00010000000000010011100011010001",	-- 7304: 	lhif	%f1, 0.000100
"00111111111111100000000000011111",	-- 7305: 	sw	%ra, [%sp + 31]
"10100111110111100000000000100000",	-- 7306: 	addi	%sp, %sp, 32
"01011000000000000000010011110011",	-- 7307: 	jal	fless.2532
"10101011110111100000000000100000",	-- 7308: 	subi	%sp, %sp, 32
"00111011110111110000000000011111",	-- 7309: 	lw	%ra, [%sp + 31]
"11001100000000100000000000000000",	-- 7310: 	lli	%r2, 0
"00101000001000100000000000010101",	-- 7311: 	bneq	%r1, %r2, bneq_else.9167
"10010011110000000000000000011001",	-- 7312: 	lf	%f0, [%sp + 25]
"10010011110000010000000000011110",	-- 7313: 	lf	%f1, [%sp + 30]
"11101100001000000000000000000000",	-- 7314: 	divf	%f0, %f1, %f0
"00111111111111100000000000011111",	-- 7315: 	sw	%ra, [%sp + 31]
"10100111110111100000000000100000",	-- 7316: 	addi	%sp, %sp, 32
"01011000000000000010101001001111",	-- 7317: 	jal	yj_fabs
"10101011110111100000000000100000",	-- 7318: 	subi	%sp, %sp, 32
"00111011110111110000000000011111",	-- 7319: 	lw	%ra, [%sp + 31]
"00111111111111100000000000011111",	-- 7320: 	sw	%ra, [%sp + 31]
"10100111110111100000000000100000",	-- 7321: 	addi	%sp, %sp, 32
"01011000000000000000010010011110",	-- 7322: 	jal	atan.2520
"10101011110111100000000000100000",	-- 7323: 	subi	%sp, %sp, 32
"00111011110111110000000000011111",	-- 7324: 	lw	%ra, [%sp + 31]
"00010100000000010000000000000000",	-- 7325: 	llif	%f1, 30.000000
"00010000000000010100000111110000",	-- 7326: 	lhif	%f1, 30.000000
"11101000000000010000000000000000",	-- 7327: 	mulf	%f0, %f0, %f1
"00010100000000010000111111011100",	-- 7328: 	llif	%f1, 3.141593
"00010000000000010100000001001001",	-- 7329: 	lhif	%f1, 3.141593
"11101100000000010000000000000000",	-- 7330: 	divf	%f0, %f0, %f1
"01010100000000000001110010100110",	-- 7331: 	j	bneq_cont.9168
	-- bneq_else.9167:
"00010100000000000000000000000000",	-- 7332: 	llif	%f0, 15.000000
"00010000000000000100000101110000",	-- 7333: 	lhif	%f0, 15.000000
	-- bneq_cont.9168:
"10110000000111100000000000011111",	-- 7334: 	sf	%f0, [%sp + 31]
"00111111111111100000000000100000",	-- 7335: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 7336: 	addi	%sp, %sp, 33
"01011000000000000010101000110010",	-- 7337: 	jal	yj_floor
"10101011110111100000000000100001",	-- 7338: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7339: 	lw	%ra, [%sp + 32]
"10010011110000010000000000011111",	-- 7340: 	lf	%f1, [%sp + 31]
"11100100001000000000000000000000",	-- 7341: 	subf	%f0, %f1, %f0
"00010100000000011001100110011010",	-- 7342: 	llif	%f1, 0.150000
"00010000000000010011111000011001",	-- 7343: 	lhif	%f1, 0.150000
"00010100000000100000000000000000",	-- 7344: 	llif	%f2, 0.500000
"00010000000000100011111100000000",	-- 7345: 	lhif	%f2, 0.500000
"10010011110000110000000000011011",	-- 7346: 	lf	%f3, [%sp + 27]
"11100100010000110001000000000000",	-- 7347: 	subf	%f2, %f2, %f3
"10110000000111100000000000100000",	-- 7348: 	sf	%f0, [%sp + 32]
"10110000001111100000000000100001",	-- 7349: 	sf	%f1, [%sp + 33]
"00001100010000000000000000000000",	-- 7350: 	movf	%f0, %f2
"00111111111111100000000000100010",	-- 7351: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 7352: 	addi	%sp, %sp, 35
"01011000000000000000010011110001",	-- 7353: 	jal	fsqr.2530
"10101011110111100000000000100011",	-- 7354: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 7355: 	lw	%ra, [%sp + 34]
"10010011110000010000000000100001",	-- 7356: 	lf	%f1, [%sp + 33]
"11100100001000000000000000000000",	-- 7357: 	subf	%f0, %f1, %f0
"00010100000000010000000000000000",	-- 7358: 	llif	%f1, 0.500000
"00010000000000010011111100000000",	-- 7359: 	lhif	%f1, 0.500000
"10010011110000100000000000100000",	-- 7360: 	lf	%f2, [%sp + 32]
"11100100001000100000100000000000",	-- 7361: 	subf	%f1, %f1, %f2
"10110000000111100000000000100010",	-- 7362: 	sf	%f0, [%sp + 34]
"00001100001000000000000000000000",	-- 7363: 	movf	%f0, %f1
"00111111111111100000000000100011",	-- 7364: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 7365: 	addi	%sp, %sp, 36
"01011000000000000000010011110001",	-- 7366: 	jal	fsqr.2530
"10101011110111100000000000100100",	-- 7367: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 7368: 	lw	%ra, [%sp + 35]
"10010011110000010000000000100010",	-- 7369: 	lf	%f1, [%sp + 34]
"11100100001000000000000000000000",	-- 7370: 	subf	%f0, %f1, %f0
"10110000000111100000000000100011",	-- 7371: 	sf	%f0, [%sp + 35]
"00111111111111100000000000100100",	-- 7372: 	sw	%ra, [%sp + 36]
"10100111110111100000000000100101",	-- 7373: 	addi	%sp, %sp, 37
"01011000000000000000010011011101",	-- 7374: 	jal	fisneg.2524
"10101011110111100000000000100101",	-- 7375: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 7376: 	lw	%ra, [%sp + 36]
"11001100000000100000000000000000",	-- 7377: 	lli	%r2, 0
"00101000001000100000000000000011",	-- 7378: 	bneq	%r1, %r2, bneq_else.9169
"10010011110000000000000000100011",	-- 7379: 	lf	%f0, [%sp + 35]
"01010100000000000001110011010111",	-- 7380: 	j	bneq_cont.9170
	-- bneq_else.9169:
"00010100000000000000000000000000",	-- 7381: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 7382: 	lhif	%f0, 0.000000
	-- bneq_cont.9170:
"11001100000000010000000000000010",	-- 7383: 	lli	%r1, 2
"00010100000000010000000000000000",	-- 7384: 	llif	%f1, 255.000000
"00010000000000010100001101111111",	-- 7385: 	lhif	%f1, 255.000000
"11101000001000000000000000000000",	-- 7386: 	mulf	%f0, %f1, %f0
"00010100000000011001100110011010",	-- 7387: 	llif	%f1, 0.300000
"00010000000000010011111010011001",	-- 7388: 	lhif	%f1, 0.300000
"11101100000000010000000000000000",	-- 7389: 	divf	%f0, %f0, %f1
"00111011110000100000000000000001",	-- 7390: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 7391: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 7392: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 7393: 	jr	%ra
	-- bneq_else.9164:
"01001111111000000000000000000000",	-- 7394: 	jr	%ra
	-- add_light.2894:
"00111011011000010000000000000010",	-- 7395: 	lw	%r1, [%r27 + 2]
"00111011011000100000000000000001",	-- 7396: 	lw	%r2, [%r27 + 1]
"10110000010111100000000000000000",	-- 7397: 	sf	%f2, [%sp + 0]
"10110000001111100000000000000001",	-- 7398: 	sf	%f1, [%sp + 1]
"10110000000111100000000000000010",	-- 7399: 	sf	%f0, [%sp + 2]
"00111100001111100000000000000011",	-- 7400: 	sw	%r1, [%sp + 3]
"00111100010111100000000000000100",	-- 7401: 	sw	%r2, [%sp + 4]
"00111111111111100000000000000101",	-- 7402: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 7403: 	addi	%sp, %sp, 6
"01011000000000000000010011010110",	-- 7404: 	jal	fispos.2522
"10101011110111100000000000000110",	-- 7405: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 7406: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000000",	-- 7407: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 7408: 	bneq	%r1, %r2, bneq_else.9173
"01010100000000000001110011111010",	-- 7409: 	j	bneq_cont.9174
	-- bneq_else.9173:
"10010011110000000000000000000010",	-- 7410: 	lf	%f0, [%sp + 2]
"00111011110000010000000000000100",	-- 7411: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000011",	-- 7412: 	lw	%r2, [%sp + 3]
"00111111111111100000000000000101",	-- 7413: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 7414: 	addi	%sp, %sp, 6
"01011000000000000000010111001110",	-- 7415: 	jal	vecaccum.2605
"10101011110111100000000000000110",	-- 7416: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 7417: 	lw	%ra, [%sp + 5]
	-- bneq_cont.9174:
"10010011110000000000000000000001",	-- 7418: 	lf	%f0, [%sp + 1]
"00111111111111100000000000000101",	-- 7419: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 7420: 	addi	%sp, %sp, 6
"01011000000000000000010011010110",	-- 7421: 	jal	fispos.2522
"10101011110111100000000000000110",	-- 7422: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 7423: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000000",	-- 7424: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 7425: 	bneq	%r1, %r2, bneq_else.9175
"01001111111000000000000000000000",	-- 7426: 	jr	%ra
	-- bneq_else.9175:
"10010011110000000000000000000001",	-- 7427: 	lf	%f0, [%sp + 1]
"00111111111111100000000000000101",	-- 7428: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 7429: 	addi	%sp, %sp, 6
"01011000000000000000010011110001",	-- 7430: 	jal	fsqr.2530
"10101011110111100000000000000110",	-- 7431: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 7432: 	lw	%ra, [%sp + 5]
"00111111111111100000000000000101",	-- 7433: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 7434: 	addi	%sp, %sp, 6
"01011000000000000000010011110001",	-- 7435: 	jal	fsqr.2530
"10101011110111100000000000000110",	-- 7436: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 7437: 	lw	%ra, [%sp + 5]
"10010011110000010000000000000000",	-- 7438: 	lf	%f1, [%sp + 0]
"11101000000000010000000000000000",	-- 7439: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000000",	-- 7440: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 7441: 	lli	%r2, 0
"00111011110000110000000000000100",	-- 7442: 	lw	%r3, [%sp + 4]
"10000100011000100001000000000000",	-- 7443: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 7444: 	lf	%f1, [%r2 + 0]
"11100000001000000000100000000000",	-- 7445: 	addf	%f1, %f1, %f0
"10000100011000010000100000000000",	-- 7446: 	add	%r1, %r3, %r1
"10110000001000010000000000000000",	-- 7447: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000001",	-- 7448: 	lli	%r1, 1
"11001100000000100000000000000001",	-- 7449: 	lli	%r2, 1
"10000100011000100001000000000000",	-- 7450: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 7451: 	lf	%f1, [%r2 + 0]
"11100000001000000000100000000000",	-- 7452: 	addf	%f1, %f1, %f0
"10000100011000010000100000000000",	-- 7453: 	add	%r1, %r3, %r1
"10110000001000010000000000000000",	-- 7454: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 7455: 	lli	%r1, 2
"11001100000000100000000000000010",	-- 7456: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 7457: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 7458: 	lf	%f1, [%r2 + 0]
"11100000001000000000000000000000",	-- 7459: 	addf	%f0, %f1, %f0
"10000100011000010000100000000000",	-- 7460: 	add	%r1, %r3, %r1
"10110000000000010000000000000000",	-- 7461: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 7462: 	jr	%ra
	-- trace_reflections.2898:
"00111011011000110000000000001000",	-- 7463: 	lw	%r3, [%r27 + 8]
"00111011011001000000000000000111",	-- 7464: 	lw	%r4, [%r27 + 7]
"00111011011001010000000000000110",	-- 7465: 	lw	%r5, [%r27 + 6]
"00111011011001100000000000000101",	-- 7466: 	lw	%r6, [%r27 + 5]
"00111011011001110000000000000100",	-- 7467: 	lw	%r7, [%r27 + 4]
"00111011011010000000000000000011",	-- 7468: 	lw	%r8, [%r27 + 3]
"00111011011010010000000000000010",	-- 7469: 	lw	%r9, [%r27 + 2]
"00111011011010100000000000000001",	-- 7470: 	lw	%r10, [%r27 + 1]
"11001100000010110000000000000000",	-- 7471: 	lli	%r11, 0
"00110001011000010000000010000001",	-- 7472: 	bgt	%r11, %r1, bgt_else.9178
"10000100100000010010000000000000",	-- 7473: 	add	%r4, %r4, %r1
"00111000100001000000000000000000",	-- 7474: 	lw	%r4, [%r4 + 0]
"00111111011111100000000000000000",	-- 7475: 	sw	%r27, [%sp + 0]
"00111100001111100000000000000001",	-- 7476: 	sw	%r1, [%sp + 1]
"10110000001111100000000000000010",	-- 7477: 	sf	%f1, [%sp + 2]
"00111101010111100000000000000011",	-- 7478: 	sw	%r10, [%sp + 3]
"00111100010111100000000000000100",	-- 7479: 	sw	%r2, [%sp + 4]
"10110000000111100000000000000101",	-- 7480: 	sf	%f0, [%sp + 5]
"00111100110111100000000000000110",	-- 7481: 	sw	%r6, [%sp + 6]
"00111100011111100000000000000111",	-- 7482: 	sw	%r3, [%sp + 7]
"00111100101111100000000000001000",	-- 7483: 	sw	%r5, [%sp + 8]
"00111100100111100000000000001001",	-- 7484: 	sw	%r4, [%sp + 9]
"00111101000111100000000000001010",	-- 7485: 	sw	%r8, [%sp + 10]
"00111101001111100000000000001011",	-- 7486: 	sw	%r9, [%sp + 11]
"00111100111111100000000000001100",	-- 7487: 	sw	%r7, [%sp + 12]
"10000100000001000000100000000000",	-- 7488: 	add	%r1, %r0, %r4
"00111111111111100000000000001101",	-- 7489: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 7490: 	addi	%sp, %sp, 14
"01011000000000000000011011000010",	-- 7491: 	jal	r_dvec.2689
"10101011110111100000000000001110",	-- 7492: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 7493: 	lw	%ra, [%sp + 13]
"00111011110110110000000000001100",	-- 7494: 	lw	%r27, [%sp + 12]
"00111100001111100000000000001101",	-- 7495: 	sw	%r1, [%sp + 13]
"00111111111111100000000000001110",	-- 7496: 	sw	%ra, [%sp + 14]
"00111011011110100000000000000000",	-- 7497: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001111",	-- 7498: 	addi	%sp, %sp, 15
"01010011010000000000000000000000",	-- 7499: 	jalr	%r26
"10101011110111100000000000001111",	-- 7500: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 7501: 	lw	%ra, [%sp + 14]
"11001100000000100000000000000000",	-- 7502: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 7503: 	bneq	%r1, %r2, bneq_else.9179
"01010100000000000001110110101000",	-- 7504: 	j	bneq_cont.9180
	-- bneq_else.9179:
"11001100000000010000000000000000",	-- 7505: 	lli	%r1, 0
"00111011110000100000000000001011",	-- 7506: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 7507: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 7508: 	lw	%r1, [%r1 + 0]
"11001100000000100000000000000100",	-- 7509: 	lli	%r2, 4
"10001100001000100000100000000000",	-- 7510: 	mul	%r1, %r1, %r2
"11001100000000100000000000000000",	-- 7511: 	lli	%r2, 0
"00111011110000110000000000001010",	-- 7512: 	lw	%r3, [%sp + 10]
"10000100011000100001000000000000",	-- 7513: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 7514: 	lw	%r2, [%r2 + 0]
"10000100001000100000100000000000",	-- 7515: 	add	%r1, %r1, %r2
"00111011110000100000000000001001",	-- 7516: 	lw	%r2, [%sp + 9]
"00111100001111100000000000001110",	-- 7517: 	sw	%r1, [%sp + 14]
"10000100000000100000100000000000",	-- 7518: 	add	%r1, %r0, %r2
"00111111111111100000000000001111",	-- 7519: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 7520: 	addi	%sp, %sp, 16
"01011000000000000000011011000000",	-- 7521: 	jal	r_surface_id.2687
"10101011110111100000000000010000",	-- 7522: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 7523: 	lw	%ra, [%sp + 15]
"00111011110000100000000000001110",	-- 7524: 	lw	%r2, [%sp + 14]
"00101000010000010000000001000011",	-- 7525: 	bneq	%r2, %r1, bneq_else.9181
"11001100000000010000000000000000",	-- 7526: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 7527: 	lli	%r2, 0
"00111011110000110000000000001000",	-- 7528: 	lw	%r3, [%sp + 8]
"10000100011000100001000000000000",	-- 7529: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 7530: 	lw	%r2, [%r2 + 0]
"00111011110110110000000000000111",	-- 7531: 	lw	%r27, [%sp + 7]
"00111111111111100000000000001111",	-- 7532: 	sw	%ra, [%sp + 15]
"00111011011110100000000000000000",	-- 7533: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010000",	-- 7534: 	addi	%sp, %sp, 16
"01010011010000000000000000000000",	-- 7535: 	jalr	%r26
"10101011110111100000000000010000",	-- 7536: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 7537: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 7538: 	lli	%r2, 0
"00101000001000100000000000110100",	-- 7539: 	bneq	%r1, %r2, bneq_else.9183
"00111011110000010000000000001101",	-- 7540: 	lw	%r1, [%sp + 13]
"00111111111111100000000000001111",	-- 7541: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 7542: 	addi	%sp, %sp, 16
"01011000000000000000011010111100",	-- 7543: 	jal	d_vec.2683
"10101011110111100000000000010000",	-- 7544: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 7545: 	lw	%ra, [%sp + 15]
"10000100000000010001000000000000",	-- 7546: 	add	%r2, %r0, %r1
"00111011110000010000000000000110",	-- 7547: 	lw	%r1, [%sp + 6]
"00111111111111100000000000001111",	-- 7548: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 7549: 	addi	%sp, %sp, 16
"01011000000000000000010110100111",	-- 7550: 	jal	veciprod.2597
"10101011110111100000000000010000",	-- 7551: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 7552: 	lw	%ra, [%sp + 15]
"00111011110000010000000000001001",	-- 7553: 	lw	%r1, [%sp + 9]
"10110000000111100000000000001111",	-- 7554: 	sf	%f0, [%sp + 15]
"00111111111111100000000000010000",	-- 7555: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 7556: 	addi	%sp, %sp, 17
"01011000000000000000011011000100",	-- 7557: 	jal	r_bright.2691
"10101011110111100000000000010001",	-- 7558: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 7559: 	lw	%ra, [%sp + 16]
"10010011110000010000000000000101",	-- 7560: 	lf	%f1, [%sp + 5]
"11101000000000010001000000000000",	-- 7561: 	mulf	%f2, %f0, %f1
"10010011110000110000000000001111",	-- 7562: 	lf	%f3, [%sp + 15]
"11101000010000110001000000000000",	-- 7563: 	mulf	%f2, %f2, %f3
"00111011110000010000000000001101",	-- 7564: 	lw	%r1, [%sp + 13]
"10110000010111100000000000010000",	-- 7565: 	sf	%f2, [%sp + 16]
"10110000000111100000000000010001",	-- 7566: 	sf	%f0, [%sp + 17]
"00111111111111100000000000010010",	-- 7567: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 7568: 	addi	%sp, %sp, 19
"01011000000000000000011010111100",	-- 7569: 	jal	d_vec.2683
"10101011110111100000000000010011",	-- 7570: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 7571: 	lw	%ra, [%sp + 18]
"10000100000000010001000000000000",	-- 7572: 	add	%r2, %r0, %r1
"00111011110000010000000000000100",	-- 7573: 	lw	%r1, [%sp + 4]
"00111111111111100000000000010010",	-- 7574: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 7575: 	addi	%sp, %sp, 19
"01011000000000000000010110100111",	-- 7576: 	jal	veciprod.2597
"10101011110111100000000000010011",	-- 7577: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 7578: 	lw	%ra, [%sp + 18]
"10010011110000010000000000010001",	-- 7579: 	lf	%f1, [%sp + 17]
"11101000001000000000100000000000",	-- 7580: 	mulf	%f1, %f1, %f0
"10010011110000000000000000010000",	-- 7581: 	lf	%f0, [%sp + 16]
"10010011110000100000000000000010",	-- 7582: 	lf	%f2, [%sp + 2]
"00111011110110110000000000000011",	-- 7583: 	lw	%r27, [%sp + 3]
"00111111111111100000000000010010",	-- 7584: 	sw	%ra, [%sp + 18]
"00111011011110100000000000000000",	-- 7585: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010011",	-- 7586: 	addi	%sp, %sp, 19
"01010011010000000000000000000000",	-- 7587: 	jalr	%r26
"10101011110111100000000000010011",	-- 7588: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 7589: 	lw	%ra, [%sp + 18]
"01010100000000000001110110100111",	-- 7590: 	j	bneq_cont.9184
	-- bneq_else.9183:
	-- bneq_cont.9184:
"01010100000000000001110110101000",	-- 7591: 	j	bneq_cont.9182
	-- bneq_else.9181:
	-- bneq_cont.9182:
	-- bneq_cont.9180:
"11001100000000010000000000000001",	-- 7592: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 7593: 	lw	%r2, [%sp + 1]
"10001000010000010000100000000000",	-- 7594: 	sub	%r1, %r2, %r1
"10010011110000000000000000000101",	-- 7595: 	lf	%f0, [%sp + 5]
"10010011110000010000000000000010",	-- 7596: 	lf	%f1, [%sp + 2]
"00111011110000100000000000000100",	-- 7597: 	lw	%r2, [%sp + 4]
"00111011110110110000000000000000",	-- 7598: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 7599: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 7600: 	jr	%r26
	-- bgt_else.9178:
"01001111111000000000000000000000",	-- 7601: 	jr	%ra
	-- trace_ray.2903:
"00111011011001000000000000010100",	-- 7602: 	lw	%r4, [%r27 + 20]
"00111011011001010000000000010011",	-- 7603: 	lw	%r5, [%r27 + 19]
"00111011011001100000000000010010",	-- 7604: 	lw	%r6, [%r27 + 18]
"00111011011001110000000000010001",	-- 7605: 	lw	%r7, [%r27 + 17]
"00111011011010000000000000010000",	-- 7606: 	lw	%r8, [%r27 + 16]
"00111011011010010000000000001111",	-- 7607: 	lw	%r9, [%r27 + 15]
"00111011011010100000000000001110",	-- 7608: 	lw	%r10, [%r27 + 14]
"00111011011010110000000000001101",	-- 7609: 	lw	%r11, [%r27 + 13]
"00111011011011000000000000001100",	-- 7610: 	lw	%r12, [%r27 + 12]
"00111011011011010000000000001011",	-- 7611: 	lw	%r13, [%r27 + 11]
"00111011011011100000000000001010",	-- 7612: 	lw	%r14, [%r27 + 10]
"00111011011011110000000000001001",	-- 7613: 	lw	%r15, [%r27 + 9]
"00111011011100000000000000001000",	-- 7614: 	lw	%r16, [%r27 + 8]
"00111011011100010000000000000111",	-- 7615: 	lw	%r17, [%r27 + 7]
"00111011011100100000000000000110",	-- 7616: 	lw	%r18, [%r27 + 6]
"00111011011100110000000000000101",	-- 7617: 	lw	%r19, [%r27 + 5]
"00111011011101000000000000000100",	-- 7618: 	lw	%r20, [%r27 + 4]
"00111011011101010000000000000011",	-- 7619: 	lw	%r21, [%r27 + 3]
"00111011011101100000000000000010",	-- 7620: 	lw	%r22, [%r27 + 2]
"00111011011101110000000000000001",	-- 7621: 	lw	%r23, [%r27 + 1]
"11001100000110000000000000000100",	-- 7622: 	lli	%r24, 4
"00110000001110000000000110101111",	-- 7623: 	bgt	%r1, %r24, bgt_else.9186
"00111111011111100000000000000000",	-- 7624: 	sw	%r27, [%sp + 0]
"10110000001111100000000000000001",	-- 7625: 	sf	%f1, [%sp + 1]
"00111100110111100000000000000010",	-- 7626: 	sw	%r6, [%sp + 2]
"00111100101111100000000000000011",	-- 7627: 	sw	%r5, [%sp + 3]
"00111101111111100000000000000100",	-- 7628: 	sw	%r15, [%sp + 4]
"00111101010111100000000000000101",	-- 7629: 	sw	%r10, [%sp + 5]
"00111110111111100000000000000110",	-- 7630: 	sw	%r23, [%sp + 6]
"00111101001111100000000000000111",	-- 7631: 	sw	%r9, [%sp + 7]
"00111101100111100000000000001000",	-- 7632: 	sw	%r12, [%sp + 8]
"00111101110111100000000000001001",	-- 7633: 	sw	%r14, [%sp + 9]
"00111100111111100000000000001010",	-- 7634: 	sw	%r7, [%sp + 10]
"00111100011111100000000000001011",	-- 7635: 	sw	%r3, [%sp + 11]
"00111110010111100000000000001100",	-- 7636: 	sw	%r18, [%sp + 12]
"00111100100111100000000000001101",	-- 7637: 	sw	%r4, [%sp + 13]
"00111110011111100000000000001110",	-- 7638: 	sw	%r19, [%sp + 14]
"00111101000111100000000000001111",	-- 7639: 	sw	%r8, [%sp + 15]
"00111110101111100000000000010000",	-- 7640: 	sw	%r21, [%sp + 16]
"00111101101111100000000000010001",	-- 7641: 	sw	%r13, [%sp + 17]
"00111110100111100000000000010010",	-- 7642: 	sw	%r20, [%sp + 18]
"00111101011111100000000000010011",	-- 7643: 	sw	%r11, [%sp + 19]
"00111110110111100000000000010100",	-- 7644: 	sw	%r22, [%sp + 20]
"10110000000111100000000000010101",	-- 7645: 	sf	%f0, [%sp + 21]
"00111110000111100000000000010110",	-- 7646: 	sw	%r16, [%sp + 22]
"00111100001111100000000000010111",	-- 7647: 	sw	%r1, [%sp + 23]
"00111100010111100000000000011000",	-- 7648: 	sw	%r2, [%sp + 24]
"00111110001111100000000000011001",	-- 7649: 	sw	%r17, [%sp + 25]
"10000100000000110000100000000000",	-- 7650: 	add	%r1, %r0, %r3
"00111111111111100000000000011010",	-- 7651: 	sw	%ra, [%sp + 26]
"10100111110111100000000000011011",	-- 7652: 	addi	%sp, %sp, 27
"01011000000000000000011010101000",	-- 7653: 	jal	p_surface_ids.2668
"10101011110111100000000000011011",	-- 7654: 	subi	%sp, %sp, 27
"00111011110111110000000000011010",	-- 7655: 	lw	%ra, [%sp + 26]
"00111011110000100000000000011000",	-- 7656: 	lw	%r2, [%sp + 24]
"00111011110110110000000000011001",	-- 7657: 	lw	%r27, [%sp + 25]
"00111100001111100000000000011010",	-- 7658: 	sw	%r1, [%sp + 26]
"10000100000000100000100000000000",	-- 7659: 	add	%r1, %r0, %r2
"00111111111111100000000000011011",	-- 7660: 	sw	%ra, [%sp + 27]
"00111011011110100000000000000000",	-- 7661: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000011100",	-- 7662: 	addi	%sp, %sp, 28
"01010011010000000000000000000000",	-- 7663: 	jalr	%r26
"10101011110111100000000000011100",	-- 7664: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 7665: 	lw	%ra, [%sp + 27]
"11001100000000100000000000000000",	-- 7666: 	lli	%r2, 0
"00101000001000100000000001000101",	-- 7667: 	bneq	%r1, %r2, bneq_else.9187
"11001100000000011111111111111111",	-- 7668: 	lli	%r1, -1
"11001000000000011111111111111111",	-- 7669: 	lhi	%r1, -1
"00111011110000100000000000010111",	-- 7670: 	lw	%r2, [%sp + 23]
"00111011110000110000000000011010",	-- 7671: 	lw	%r3, [%sp + 26]
"10000100011000100001100000000000",	-- 7672: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 7673: 	sw	%r1, [%r3 + 0]
"11001100000000010000000000000000",	-- 7674: 	lli	%r1, 0
"00101000010000010000000000000010",	-- 7675: 	bneq	%r2, %r1, bneq_else.9188
"01001111111000000000000000000000",	-- 7676: 	jr	%ra
	-- bneq_else.9188:
"00111011110000010000000000011000",	-- 7677: 	lw	%r1, [%sp + 24]
"00111011110000100000000000010110",	-- 7678: 	lw	%r2, [%sp + 22]
"00111111111111100000000000011011",	-- 7679: 	sw	%ra, [%sp + 27]
"10100111110111100000000000011100",	-- 7680: 	addi	%sp, %sp, 28
"01011000000000000000010110100111",	-- 7681: 	jal	veciprod.2597
"10101011110111100000000000011100",	-- 7682: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 7683: 	lw	%ra, [%sp + 27]
"00111111111111100000000000011011",	-- 7684: 	sw	%ra, [%sp + 27]
"10100111110111100000000000011100",	-- 7685: 	addi	%sp, %sp, 28
"01011000000000000010101001010001",	-- 7686: 	jal	yj_fneg
"10101011110111100000000000011100",	-- 7687: 	subi	%sp, %sp, 28
"00111011110111110000000000011011",	-- 7688: 	lw	%ra, [%sp + 27]
"10110000000111100000000000011011",	-- 7689: 	sf	%f0, [%sp + 27]
"00111111111111100000000000011100",	-- 7690: 	sw	%ra, [%sp + 28]
"10100111110111100000000000011101",	-- 7691: 	addi	%sp, %sp, 29
"01011000000000000000010011010110",	-- 7692: 	jal	fispos.2522
"10101011110111100000000000011101",	-- 7693: 	subi	%sp, %sp, 29
"00111011110111110000000000011100",	-- 7694: 	lw	%ra, [%sp + 28]
"11001100000000100000000000000000",	-- 7695: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 7696: 	bneq	%r1, %r2, bneq_else.9190
"01001111111000000000000000000000",	-- 7697: 	jr	%ra
	-- bneq_else.9190:
"10010011110000000000000000011011",	-- 7698: 	lf	%f0, [%sp + 27]
"00111111111111100000000000011100",	-- 7699: 	sw	%ra, [%sp + 28]
"10100111110111100000000000011101",	-- 7700: 	addi	%sp, %sp, 29
"01011000000000000000010011110001",	-- 7701: 	jal	fsqr.2530
"10101011110111100000000000011101",	-- 7702: 	subi	%sp, %sp, 29
"00111011110111110000000000011100",	-- 7703: 	lw	%ra, [%sp + 28]
"10010011110000010000000000011011",	-- 7704: 	lf	%f1, [%sp + 27]
"11101000000000010000000000000000",	-- 7705: 	mulf	%f0, %f0, %f1
"10010011110000010000000000010101",	-- 7706: 	lf	%f1, [%sp + 21]
"11101000000000010000000000000000",	-- 7707: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000000",	-- 7708: 	lli	%r1, 0
"00111011110000100000000000010100",	-- 7709: 	lw	%r2, [%sp + 20]
"10000100010000010000100000000000",	-- 7710: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 7711: 	lf	%f1, [%r1 + 0]
"11101000000000010000000000000000",	-- 7712: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000000",	-- 7713: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 7714: 	lli	%r2, 0
"00111011110000110000000000010011",	-- 7715: 	lw	%r3, [%sp + 19]
"10000100011000100001000000000000",	-- 7716: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 7717: 	lf	%f1, [%r2 + 0]
"11100000001000000000100000000000",	-- 7718: 	addf	%f1, %f1, %f0
"10000100011000010000100000000000",	-- 7719: 	add	%r1, %r3, %r1
"10110000001000010000000000000000",	-- 7720: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000001",	-- 7721: 	lli	%r1, 1
"11001100000000100000000000000001",	-- 7722: 	lli	%r2, 1
"10000100011000100001000000000000",	-- 7723: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 7724: 	lf	%f1, [%r2 + 0]
"11100000001000000000100000000000",	-- 7725: 	addf	%f1, %f1, %f0
"10000100011000010000100000000000",	-- 7726: 	add	%r1, %r3, %r1
"10110000001000010000000000000000",	-- 7727: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 7728: 	lli	%r1, 2
"11001100000000100000000000000010",	-- 7729: 	lli	%r2, 2
"10000100011000100001000000000000",	-- 7730: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 7731: 	lf	%f1, [%r2 + 0]
"11100000001000000000000000000000",	-- 7732: 	addf	%f0, %f1, %f0
"10000100011000010000100000000000",	-- 7733: 	add	%r1, %r3, %r1
"10110000000000010000000000000000",	-- 7734: 	sf	%f0, [%r1 + 0]
"01001111111000000000000000000000",	-- 7735: 	jr	%ra
	-- bneq_else.9187:
"11001100000000010000000000000000",	-- 7736: 	lli	%r1, 0
"00111011110000100000000000010010",	-- 7737: 	lw	%r2, [%sp + 18]
"10000100010000010000100000000000",	-- 7738: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 7739: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000010001",	-- 7740: 	lw	%r2, [%sp + 17]
"10000100010000010001000000000000",	-- 7741: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 7742: 	lw	%r2, [%r2 + 0]
"00111100001111100000000000011100",	-- 7743: 	sw	%r1, [%sp + 28]
"00111100010111100000000000011101",	-- 7744: 	sw	%r2, [%sp + 29]
"10000100000000100000100000000000",	-- 7745: 	add	%r1, %r0, %r2
"00111111111111100000000000011110",	-- 7746: 	sw	%ra, [%sp + 30]
"10100111110111100000000000011111",	-- 7747: 	addi	%sp, %sp, 31
"01011000000000000000011001010100",	-- 7748: 	jal	o_reflectiontype.2626
"10101011110111100000000000011111",	-- 7749: 	subi	%sp, %sp, 31
"00111011110111110000000000011110",	-- 7750: 	lw	%ra, [%sp + 30]
"00111011110000100000000000011101",	-- 7751: 	lw	%r2, [%sp + 29]
"00111100001111100000000000011110",	-- 7752: 	sw	%r1, [%sp + 30]
"10000100000000100000100000000000",	-- 7753: 	add	%r1, %r0, %r2
"00111111111111100000000000011111",	-- 7754: 	sw	%ra, [%sp + 31]
"10100111110111100000000000100000",	-- 7755: 	addi	%sp, %sp, 32
"01011000000000000000011001111010",	-- 7756: 	jal	o_diffuse.2646
"10101011110111100000000000100000",	-- 7757: 	subi	%sp, %sp, 32
"00111011110111110000000000011111",	-- 7758: 	lw	%ra, [%sp + 31]
"10010011110000010000000000010101",	-- 7759: 	lf	%f1, [%sp + 21]
"11101000000000010000000000000000",	-- 7760: 	mulf	%f0, %f0, %f1
"00111011110000010000000000011101",	-- 7761: 	lw	%r1, [%sp + 29]
"00111011110000100000000000011000",	-- 7762: 	lw	%r2, [%sp + 24]
"00111011110110110000000000010000",	-- 7763: 	lw	%r27, [%sp + 16]
"10110000000111100000000000011111",	-- 7764: 	sf	%f0, [%sp + 31]
"00111111111111100000000000100000",	-- 7765: 	sw	%ra, [%sp + 32]
"00111011011110100000000000000000",	-- 7766: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100001",	-- 7767: 	addi	%sp, %sp, 33
"01010011010000000000000000000000",	-- 7768: 	jalr	%r26
"10101011110111100000000000100001",	-- 7769: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7770: 	lw	%ra, [%sp + 32]
"00111011110000010000000000001111",	-- 7771: 	lw	%r1, [%sp + 15]
"00111011110000100000000000001110",	-- 7772: 	lw	%r2, [%sp + 14]
"00111111111111100000000000100000",	-- 7773: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 7774: 	addi	%sp, %sp, 33
"01011000000000000000010100111101",	-- 7775: 	jal	veccpy.2586
"10101011110111100000000000100001",	-- 7776: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7777: 	lw	%ra, [%sp + 32]
"00111011110000010000000000011101",	-- 7778: 	lw	%r1, [%sp + 29]
"00111011110000100000000000001110",	-- 7779: 	lw	%r2, [%sp + 14]
"00111011110110110000000000001101",	-- 7780: 	lw	%r27, [%sp + 13]
"00111111111111100000000000100000",	-- 7781: 	sw	%ra, [%sp + 32]
"00111011011110100000000000000000",	-- 7782: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100001",	-- 7783: 	addi	%sp, %sp, 33
"01010011010000000000000000000000",	-- 7784: 	jalr	%r26
"10101011110111100000000000100001",	-- 7785: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7786: 	lw	%ra, [%sp + 32]
"11001100000000010000000000000100",	-- 7787: 	lli	%r1, 4
"00111011110000100000000000011100",	-- 7788: 	lw	%r2, [%sp + 28]
"10001100010000010000100000000000",	-- 7789: 	mul	%r1, %r2, %r1
"11001100000000100000000000000000",	-- 7790: 	lli	%r2, 0
"00111011110000110000000000001100",	-- 7791: 	lw	%r3, [%sp + 12]
"10000100011000100001000000000000",	-- 7792: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 7793: 	lw	%r2, [%r2 + 0]
"10000100001000100000100000000000",	-- 7794: 	add	%r1, %r1, %r2
"00111011110000100000000000010111",	-- 7795: 	lw	%r2, [%sp + 23]
"00111011110000110000000000011010",	-- 7796: 	lw	%r3, [%sp + 26]
"10000100011000100010000000000000",	-- 7797: 	add	%r4, %r3, %r2
"00111100001001000000000000000000",	-- 7798: 	sw	%r1, [%r4 + 0]
"00111011110000010000000000001011",	-- 7799: 	lw	%r1, [%sp + 11]
"00111111111111100000000000100000",	-- 7800: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 7801: 	addi	%sp, %sp, 33
"01011000000000000000011010100110",	-- 7802: 	jal	p_intersection_points.2666
"10101011110111100000000000100001",	-- 7803: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7804: 	lw	%ra, [%sp + 32]
"00111011110000100000000000010111",	-- 7805: 	lw	%r2, [%sp + 23]
"10000100001000100000100000000000",	-- 7806: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 7807: 	lw	%r1, [%r1 + 0]
"00111011110000110000000000001110",	-- 7808: 	lw	%r3, [%sp + 14]
"10000100000000110001000000000000",	-- 7809: 	add	%r2, %r0, %r3
"00111111111111100000000000100000",	-- 7810: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 7811: 	addi	%sp, %sp, 33
"01011000000000000000010100111101",	-- 7812: 	jal	veccpy.2586
"10101011110111100000000000100001",	-- 7813: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7814: 	lw	%ra, [%sp + 32]
"00111011110000010000000000001011",	-- 7815: 	lw	%r1, [%sp + 11]
"00111111111111100000000000100000",	-- 7816: 	sw	%ra, [%sp + 32]
"10100111110111100000000000100001",	-- 7817: 	addi	%sp, %sp, 33
"01011000000000000000011010101010",	-- 7818: 	jal	p_calc_diffuse.2670
"10101011110111100000000000100001",	-- 7819: 	subi	%sp, %sp, 33
"00111011110111110000000000100000",	-- 7820: 	lw	%ra, [%sp + 32]
"00111011110000100000000000011101",	-- 7821: 	lw	%r2, [%sp + 29]
"00111100001111100000000000100000",	-- 7822: 	sw	%r1, [%sp + 32]
"10000100000000100000100000000000",	-- 7823: 	add	%r1, %r0, %r2
"00111111111111100000000000100001",	-- 7824: 	sw	%ra, [%sp + 33]
"10100111110111100000000000100010",	-- 7825: 	addi	%sp, %sp, 34
"01011000000000000000011001111010",	-- 7826: 	jal	o_diffuse.2646
"10101011110111100000000000100010",	-- 7827: 	subi	%sp, %sp, 34
"00111011110111110000000000100001",	-- 7828: 	lw	%ra, [%sp + 33]
"00010100000000010000000000000000",	-- 7829: 	llif	%f1, 0.500000
"00010000000000010011111100000000",	-- 7830: 	lhif	%f1, 0.500000
"00111111111111100000000000100001",	-- 7831: 	sw	%ra, [%sp + 33]
"10100111110111100000000000100010",	-- 7832: 	addi	%sp, %sp, 34
"01011000000000000000010011110011",	-- 7833: 	jal	fless.2532
"10101011110111100000000000100010",	-- 7834: 	subi	%sp, %sp, 34
"00111011110111110000000000100001",	-- 7835: 	lw	%ra, [%sp + 33]
"11001100000000100000000000000000",	-- 7836: 	lli	%r2, 0
"00101000001000100000000000110111",	-- 7837: 	bneq	%r1, %r2, bneq_else.9193
"11001100000000010000000000000001",	-- 7838: 	lli	%r1, 1
"00111011110000100000000000010111",	-- 7839: 	lw	%r2, [%sp + 23]
"00111011110000110000000000100000",	-- 7840: 	lw	%r3, [%sp + 32]
"10000100011000100001100000000000",	-- 7841: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 7842: 	sw	%r1, [%r3 + 0]
"00111011110000010000000000001011",	-- 7843: 	lw	%r1, [%sp + 11]
"00111111111111100000000000100001",	-- 7844: 	sw	%ra, [%sp + 33]
"10100111110111100000000000100010",	-- 7845: 	addi	%sp, %sp, 34
"01011000000000000000011010101100",	-- 7846: 	jal	p_energy.2672
"10101011110111100000000000100010",	-- 7847: 	subi	%sp, %sp, 34
"00111011110111110000000000100001",	-- 7848: 	lw	%ra, [%sp + 33]
"00111011110000100000000000010111",	-- 7849: 	lw	%r2, [%sp + 23]
"10000100001000100001100000000000",	-- 7850: 	add	%r3, %r1, %r2
"00111000011000110000000000000000",	-- 7851: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000001010",	-- 7852: 	lw	%r4, [%sp + 10]
"00111100001111100000000000100001",	-- 7853: 	sw	%r1, [%sp + 33]
"10000100000001000001000000000000",	-- 7854: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 7855: 	add	%r1, %r0, %r3
"00111111111111100000000000100010",	-- 7856: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 7857: 	addi	%sp, %sp, 35
"01011000000000000000010100111101",	-- 7858: 	jal	veccpy.2586
"10101011110111100000000000100011",	-- 7859: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 7860: 	lw	%ra, [%sp + 34]
"00111011110000010000000000010111",	-- 7861: 	lw	%r1, [%sp + 23]
"00111011110000100000000000100001",	-- 7862: 	lw	%r2, [%sp + 33]
"10000100010000010001000000000000",	-- 7863: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 7864: 	lw	%r2, [%r2 + 0]
"00010100000000001111101111001110",	-- 7865: 	llif	%f0, 0.003906
"00010000000000000011101101111111",	-- 7866: 	lhif	%f0, 0.003906
"10010011110000010000000000011111",	-- 7867: 	lf	%f1, [%sp + 31]
"11101000000000010000000000000000",	-- 7868: 	mulf	%f0, %f0, %f1
"10000100000000100000100000000000",	-- 7869: 	add	%r1, %r0, %r2
"00111111111111100000000000100010",	-- 7870: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 7871: 	addi	%sp, %sp, 35
"01011000000000000000011000001111",	-- 7872: 	jal	vecscale.2615
"10101011110111100000000000100011",	-- 7873: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 7874: 	lw	%ra, [%sp + 34]
"00111011110000010000000000001011",	-- 7875: 	lw	%r1, [%sp + 11]
"00111111111111100000000000100010",	-- 7876: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 7877: 	addi	%sp, %sp, 35
"01011000000000000000011010111010",	-- 7878: 	jal	p_nvectors.2681
"10101011110111100000000000100011",	-- 7879: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 7880: 	lw	%ra, [%sp + 34]
"00111011110000100000000000010111",	-- 7881: 	lw	%r2, [%sp + 23]
"10000100001000100000100000000000",	-- 7882: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 7883: 	lw	%r1, [%r1 + 0]
"00111011110000110000000000001001",	-- 7884: 	lw	%r3, [%sp + 9]
"10000100000000110001000000000000",	-- 7885: 	add	%r2, %r0, %r3
"00111111111111100000000000100010",	-- 7886: 	sw	%ra, [%sp + 34]
"10100111110111100000000000100011",	-- 7887: 	addi	%sp, %sp, 35
"01011000000000000000010100111101",	-- 7888: 	jal	veccpy.2586
"10101011110111100000000000100011",	-- 7889: 	subi	%sp, %sp, 35
"00111011110111110000000000100010",	-- 7890: 	lw	%ra, [%sp + 34]
"01010100000000000001111011011001",	-- 7891: 	j	bneq_cont.9194
	-- bneq_else.9193:
"11001100000000010000000000000000",	-- 7892: 	lli	%r1, 0
"00111011110000100000000000010111",	-- 7893: 	lw	%r2, [%sp + 23]
"00111011110000110000000000100000",	-- 7894: 	lw	%r3, [%sp + 32]
"10000100011000100001100000000000",	-- 7895: 	add	%r3, %r3, %r2
"00111100001000110000000000000000",	-- 7896: 	sw	%r1, [%r3 + 0]
	-- bneq_cont.9194:
"00010100000000000000000000000000",	-- 7897: 	llif	%f0, -2.000000
"00010000000000001100000000000000",	-- 7898: 	lhif	%f0, -2.000000
"00111011110000010000000000011000",	-- 7899: 	lw	%r1, [%sp + 24]
"00111011110000100000000000001001",	-- 7900: 	lw	%r2, [%sp + 9]
"10110000000111100000000000100010",	-- 7901: 	sf	%f0, [%sp + 34]
"00111111111111100000000000100011",	-- 7902: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 7903: 	addi	%sp, %sp, 36
"01011000000000000000010110100111",	-- 7904: 	jal	veciprod.2597
"10101011110111100000000000100100",	-- 7905: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 7906: 	lw	%ra, [%sp + 35]
"10010011110000010000000000100010",	-- 7907: 	lf	%f1, [%sp + 34]
"11101000001000000000000000000000",	-- 7908: 	mulf	%f0, %f1, %f0
"00111011110000010000000000011000",	-- 7909: 	lw	%r1, [%sp + 24]
"00111011110000100000000000001001",	-- 7910: 	lw	%r2, [%sp + 9]
"00111111111111100000000000100011",	-- 7911: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 7912: 	addi	%sp, %sp, 36
"01011000000000000000010111001110",	-- 7913: 	jal	vecaccum.2605
"10101011110111100000000000100100",	-- 7914: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 7915: 	lw	%ra, [%sp + 35]
"00111011110000010000000000011101",	-- 7916: 	lw	%r1, [%sp + 29]
"00111111111111100000000000100011",	-- 7917: 	sw	%ra, [%sp + 35]
"10100111110111100000000000100100",	-- 7918: 	addi	%sp, %sp, 36
"01011000000000000000011001111111",	-- 7919: 	jal	o_hilight.2648
"10101011110111100000000000100100",	-- 7920: 	subi	%sp, %sp, 36
"00111011110111110000000000100011",	-- 7921: 	lw	%ra, [%sp + 35]
"10010011110000010000000000010101",	-- 7922: 	lf	%f1, [%sp + 21]
"11101000001000000000000000000000",	-- 7923: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 7924: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 7925: 	lli	%r2, 0
"00111011110000110000000000001000",	-- 7926: 	lw	%r3, [%sp + 8]
"10000100011000100001000000000000",	-- 7927: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 7928: 	lw	%r2, [%r2 + 0]
"00111011110110110000000000000111",	-- 7929: 	lw	%r27, [%sp + 7]
"10110000000111100000000000100011",	-- 7930: 	sf	%f0, [%sp + 35]
"00111111111111100000000000100100",	-- 7931: 	sw	%ra, [%sp + 36]
"00111011011110100000000000000000",	-- 7932: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100101",	-- 7933: 	addi	%sp, %sp, 37
"01010011010000000000000000000000",	-- 7934: 	jalr	%r26
"10101011110111100000000000100101",	-- 7935: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 7936: 	lw	%ra, [%sp + 36]
"11001100000000100000000000000000",	-- 7937: 	lli	%r2, 0
"00101000001000100000000000100111",	-- 7938: 	bneq	%r1, %r2, bneq_else.9195
"00111011110000010000000000001001",	-- 7939: 	lw	%r1, [%sp + 9]
"00111011110000100000000000010110",	-- 7940: 	lw	%r2, [%sp + 22]
"00111111111111100000000000100100",	-- 7941: 	sw	%ra, [%sp + 36]
"10100111110111100000000000100101",	-- 7942: 	addi	%sp, %sp, 37
"01011000000000000000010110100111",	-- 7943: 	jal	veciprod.2597
"10101011110111100000000000100101",	-- 7944: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 7945: 	lw	%ra, [%sp + 36]
"00111111111111100000000000100100",	-- 7946: 	sw	%ra, [%sp + 36]
"10100111110111100000000000100101",	-- 7947: 	addi	%sp, %sp, 37
"01011000000000000010101001010001",	-- 7948: 	jal	yj_fneg
"10101011110111100000000000100101",	-- 7949: 	subi	%sp, %sp, 37
"00111011110111110000000000100100",	-- 7950: 	lw	%ra, [%sp + 36]
"10010011110000010000000000011111",	-- 7951: 	lf	%f1, [%sp + 31]
"11101000000000010000000000000000",	-- 7952: 	mulf	%f0, %f0, %f1
"00111011110000010000000000011000",	-- 7953: 	lw	%r1, [%sp + 24]
"00111011110000100000000000010110",	-- 7954: 	lw	%r2, [%sp + 22]
"10110000000111100000000000100100",	-- 7955: 	sf	%f0, [%sp + 36]
"00111111111111100000000000100101",	-- 7956: 	sw	%ra, [%sp + 37]
"10100111110111100000000000100110",	-- 7957: 	addi	%sp, %sp, 38
"01011000000000000000010110100111",	-- 7958: 	jal	veciprod.2597
"10101011110111100000000000100110",	-- 7959: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 7960: 	lw	%ra, [%sp + 37]
"00111111111111100000000000100101",	-- 7961: 	sw	%ra, [%sp + 37]
"10100111110111100000000000100110",	-- 7962: 	addi	%sp, %sp, 38
"01011000000000000010101001010001",	-- 7963: 	jal	yj_fneg
"10101011110111100000000000100110",	-- 7964: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 7965: 	lw	%ra, [%sp + 37]
"00001100000000010000000000000000",	-- 7966: 	movf	%f1, %f0
"10010011110000000000000000100100",	-- 7967: 	lf	%f0, [%sp + 36]
"10010011110000100000000000100011",	-- 7968: 	lf	%f2, [%sp + 35]
"00111011110110110000000000000110",	-- 7969: 	lw	%r27, [%sp + 6]
"00111111111111100000000000100101",	-- 7970: 	sw	%ra, [%sp + 37]
"00111011011110100000000000000000",	-- 7971: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100110",	-- 7972: 	addi	%sp, %sp, 38
"01010011010000000000000000000000",	-- 7973: 	jalr	%r26
"10101011110111100000000000100110",	-- 7974: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 7975: 	lw	%ra, [%sp + 37]
"01010100000000000001111100101001",	-- 7976: 	j	bneq_cont.9196
	-- bneq_else.9195:
	-- bneq_cont.9196:
"00111011110000010000000000001110",	-- 7977: 	lw	%r1, [%sp + 14]
"00111011110110110000000000000101",	-- 7978: 	lw	%r27, [%sp + 5]
"00111111111111100000000000100101",	-- 7979: 	sw	%ra, [%sp + 37]
"00111011011110100000000000000000",	-- 7980: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100110",	-- 7981: 	addi	%sp, %sp, 38
"01010011010000000000000000000000",	-- 7982: 	jalr	%r26
"10101011110111100000000000100110",	-- 7983: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 7984: 	lw	%ra, [%sp + 37]
"11001100000000010000000000000000",	-- 7985: 	lli	%r1, 0
"00111011110000100000000000000100",	-- 7986: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 7987: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 7988: 	lw	%r1, [%r1 + 0]
"11001100000000100000000000000001",	-- 7989: 	lli	%r2, 1
"10001000001000100000100000000000",	-- 7990: 	sub	%r1, %r1, %r2
"10010011110000000000000000011111",	-- 7991: 	lf	%f0, [%sp + 31]
"10010011110000010000000000100011",	-- 7992: 	lf	%f1, [%sp + 35]
"00111011110000100000000000011000",	-- 7993: 	lw	%r2, [%sp + 24]
"00111011110110110000000000000011",	-- 7994: 	lw	%r27, [%sp + 3]
"00111111111111100000000000100101",	-- 7995: 	sw	%ra, [%sp + 37]
"00111011011110100000000000000000",	-- 7996: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000100110",	-- 7997: 	addi	%sp, %sp, 38
"01010011010000000000000000000000",	-- 7998: 	jalr	%r26
"10101011110111100000000000100110",	-- 7999: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 8000: 	lw	%ra, [%sp + 37]
"00010100000000001100110011001101",	-- 8001: 	llif	%f0, 0.100000
"00010000000000000011110111001100",	-- 8002: 	lhif	%f0, 0.100000
"10010011110000010000000000010101",	-- 8003: 	lf	%f1, [%sp + 21]
"00111111111111100000000000100101",	-- 8004: 	sw	%ra, [%sp + 37]
"10100111110111100000000000100110",	-- 8005: 	addi	%sp, %sp, 38
"01011000000000000000010011110011",	-- 8006: 	jal	fless.2532
"10101011110111100000000000100110",	-- 8007: 	subi	%sp, %sp, 38
"00111011110111110000000000100101",	-- 8008: 	lw	%ra, [%sp + 37]
"11001100000000100000000000000000",	-- 8009: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 8010: 	bneq	%r1, %r2, bneq_else.9197
"01001111111000000000000000000000",	-- 8011: 	jr	%ra
	-- bneq_else.9197:
"11001100000000010000000000000100",	-- 8012: 	lli	%r1, 4
"00111011110000100000000000010111",	-- 8013: 	lw	%r2, [%sp + 23]
"00110000001000100000000000000010",	-- 8014: 	bgt	%r1, %r2, bgt_else.9199
"01010100000000000001111101010111",	-- 8015: 	j	bgt_cont.9200
	-- bgt_else.9199:
"11001100000000010000000000000001",	-- 8016: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 8017: 	add	%r1, %r2, %r1
"11001100000000111111111111111111",	-- 8018: 	lli	%r3, -1
"11001000000000111111111111111111",	-- 8019: 	lhi	%r3, -1
"00111011110001000000000000011010",	-- 8020: 	lw	%r4, [%sp + 26]
"10000100100000010000100000000000",	-- 8021: 	add	%r1, %r4, %r1
"00111100011000010000000000000000",	-- 8022: 	sw	%r3, [%r1 + 0]
	-- bgt_cont.9200:
"11001100000000010000000000000010",	-- 8023: 	lli	%r1, 2
"00111011110000110000000000011110",	-- 8024: 	lw	%r3, [%sp + 30]
"00101000011000010000000000011100",	-- 8025: 	bneq	%r3, %r1, bneq_else.9201
"00010100000000000000000000000000",	-- 8026: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 8027: 	lhif	%f0, 1.000000
"00111011110000010000000000011101",	-- 8028: 	lw	%r1, [%sp + 29]
"10110000000111100000000000100101",	-- 8029: 	sf	%f0, [%sp + 37]
"00111111111111100000000000100110",	-- 8030: 	sw	%ra, [%sp + 38]
"10100111110111100000000000100111",	-- 8031: 	addi	%sp, %sp, 39
"01011000000000000000011001111010",	-- 8032: 	jal	o_diffuse.2646
"10101011110111100000000000100111",	-- 8033: 	subi	%sp, %sp, 39
"00111011110111110000000000100110",	-- 8034: 	lw	%ra, [%sp + 38]
"10010011110000010000000000100101",	-- 8035: 	lf	%f1, [%sp + 37]
"11100100001000000000000000000000",	-- 8036: 	subf	%f0, %f1, %f0
"10010011110000010000000000010101",	-- 8037: 	lf	%f1, [%sp + 21]
"11101000001000000000000000000000",	-- 8038: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000001",	-- 8039: 	lli	%r1, 1
"00111011110000100000000000010111",	-- 8040: 	lw	%r2, [%sp + 23]
"10000100010000010000100000000000",	-- 8041: 	add	%r1, %r2, %r1
"11001100000000100000000000000000",	-- 8042: 	lli	%r2, 0
"00111011110000110000000000000010",	-- 8043: 	lw	%r3, [%sp + 2]
"10000100011000100001000000000000",	-- 8044: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 8045: 	lf	%f1, [%r2 + 0]
"10010011110000100000000000000001",	-- 8046: 	lf	%f2, [%sp + 1]
"11100000010000010000100000000000",	-- 8047: 	addf	%f1, %f2, %f1
"00111011110000100000000000011000",	-- 8048: 	lw	%r2, [%sp + 24]
"00111011110000110000000000001011",	-- 8049: 	lw	%r3, [%sp + 11]
"00111011110110110000000000000000",	-- 8050: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 8051: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8052: 	jr	%r26
	-- bneq_else.9201:
"01001111111000000000000000000000",	-- 8053: 	jr	%ra
	-- bgt_else.9186:
"01001111111000000000000000000000",	-- 8054: 	jr	%ra
	-- trace_diffuse_ray.2909:
"00111011011000100000000000001100",	-- 8055: 	lw	%r2, [%r27 + 12]
"00111011011000110000000000001011",	-- 8056: 	lw	%r3, [%r27 + 11]
"00111011011001000000000000001010",	-- 8057: 	lw	%r4, [%r27 + 10]
"00111011011001010000000000001001",	-- 8058: 	lw	%r5, [%r27 + 9]
"00111011011001100000000000001000",	-- 8059: 	lw	%r6, [%r27 + 8]
"00111011011001110000000000000111",	-- 8060: 	lw	%r7, [%r27 + 7]
"00111011011010000000000000000110",	-- 8061: 	lw	%r8, [%r27 + 6]
"00111011011010010000000000000101",	-- 8062: 	lw	%r9, [%r27 + 5]
"00111011011010100000000000000100",	-- 8063: 	lw	%r10, [%r27 + 4]
"00111011011010110000000000000011",	-- 8064: 	lw	%r11, [%r27 + 3]
"00111011011011000000000000000010",	-- 8065: 	lw	%r12, [%r27 + 2]
"00111011011011010000000000000001",	-- 8066: 	lw	%r13, [%r27 + 1]
"00111100011111100000000000000000",	-- 8067: 	sw	%r3, [%sp + 0]
"00111101101111100000000000000001",	-- 8068: 	sw	%r13, [%sp + 1]
"10110000000111100000000000000010",	-- 8069: 	sf	%f0, [%sp + 2]
"00111101000111100000000000000011",	-- 8070: 	sw	%r8, [%sp + 3]
"00111100111111100000000000000100",	-- 8071: 	sw	%r7, [%sp + 4]
"00111100100111100000000000000101",	-- 8072: 	sw	%r4, [%sp + 5]
"00111100101111100000000000000110",	-- 8073: 	sw	%r5, [%sp + 6]
"00111101010111100000000000000111",	-- 8074: 	sw	%r10, [%sp + 7]
"00111100010111100000000000001000",	-- 8075: 	sw	%r2, [%sp + 8]
"00111101100111100000000000001001",	-- 8076: 	sw	%r12, [%sp + 9]
"00111100001111100000000000001010",	-- 8077: 	sw	%r1, [%sp + 10]
"00111100110111100000000000001011",	-- 8078: 	sw	%r6, [%sp + 11]
"00111101011111100000000000001100",	-- 8079: 	sw	%r11, [%sp + 12]
"10000100000010011101100000000000",	-- 8080: 	add	%r27, %r0, %r9
"00111111111111100000000000001101",	-- 8081: 	sw	%ra, [%sp + 13]
"00111011011110100000000000000000",	-- 8082: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001110",	-- 8083: 	addi	%sp, %sp, 14
"01010011010000000000000000000000",	-- 8084: 	jalr	%r26
"10101011110111100000000000001110",	-- 8085: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 8086: 	lw	%ra, [%sp + 13]
"11001100000000100000000000000000",	-- 8087: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 8088: 	bneq	%r1, %r2, bneq_else.9204
"01001111111000000000000000000000",	-- 8089: 	jr	%ra
	-- bneq_else.9204:
"11001100000000010000000000000000",	-- 8090: 	lli	%r1, 0
"00111011110000100000000000001100",	-- 8091: 	lw	%r2, [%sp + 12]
"10000100010000010000100000000000",	-- 8092: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8093: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000001011",	-- 8094: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 8095: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8096: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000001010",	-- 8097: 	lw	%r2, [%sp + 10]
"00111100001111100000000000001101",	-- 8098: 	sw	%r1, [%sp + 13]
"10000100000000100000100000000000",	-- 8099: 	add	%r1, %r0, %r2
"00111111111111100000000000001110",	-- 8100: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 8101: 	addi	%sp, %sp, 15
"01011000000000000000011010111100",	-- 8102: 	jal	d_vec.2683
"10101011110111100000000000001111",	-- 8103: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 8104: 	lw	%ra, [%sp + 14]
"10000100000000010001000000000000",	-- 8105: 	add	%r2, %r0, %r1
"00111011110000010000000000001101",	-- 8106: 	lw	%r1, [%sp + 13]
"00111011110110110000000000001001",	-- 8107: 	lw	%r27, [%sp + 9]
"00111111111111100000000000001110",	-- 8108: 	sw	%ra, [%sp + 14]
"00111011011110100000000000000000",	-- 8109: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001111",	-- 8110: 	addi	%sp, %sp, 15
"01010011010000000000000000000000",	-- 8111: 	jalr	%r26
"10101011110111100000000000001111",	-- 8112: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 8113: 	lw	%ra, [%sp + 14]
"00111011110000010000000000001101",	-- 8114: 	lw	%r1, [%sp + 13]
"00111011110000100000000000000111",	-- 8115: 	lw	%r2, [%sp + 7]
"00111011110110110000000000001000",	-- 8116: 	lw	%r27, [%sp + 8]
"00111111111111100000000000001110",	-- 8117: 	sw	%ra, [%sp + 14]
"00111011011110100000000000000000",	-- 8118: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001111",	-- 8119: 	addi	%sp, %sp, 15
"01010011010000000000000000000000",	-- 8120: 	jalr	%r26
"10101011110111100000000000001111",	-- 8121: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 8122: 	lw	%ra, [%sp + 14]
"11001100000000010000000000000000",	-- 8123: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 8124: 	lli	%r2, 0
"00111011110000110000000000000110",	-- 8125: 	lw	%r3, [%sp + 6]
"10000100011000100001000000000000",	-- 8126: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 8127: 	lw	%r2, [%r2 + 0]
"00111011110110110000000000000101",	-- 8128: 	lw	%r27, [%sp + 5]
"00111111111111100000000000001110",	-- 8129: 	sw	%ra, [%sp + 14]
"00111011011110100000000000000000",	-- 8130: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001111",	-- 8131: 	addi	%sp, %sp, 15
"01010011010000000000000000000000",	-- 8132: 	jalr	%r26
"10101011110111100000000000001111",	-- 8133: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 8134: 	lw	%ra, [%sp + 14]
"11001100000000100000000000000000",	-- 8135: 	lli	%r2, 0
"00101000001000100000000000100111",	-- 8136: 	bneq	%r1, %r2, bneq_else.9206
"00111011110000010000000000000100",	-- 8137: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000011",	-- 8138: 	lw	%r2, [%sp + 3]
"00111111111111100000000000001110",	-- 8139: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 8140: 	addi	%sp, %sp, 15
"01011000000000000000010110100111",	-- 8141: 	jal	veciprod.2597
"10101011110111100000000000001111",	-- 8142: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 8143: 	lw	%ra, [%sp + 14]
"00111111111111100000000000001110",	-- 8144: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 8145: 	addi	%sp, %sp, 15
"01011000000000000010101001010001",	-- 8146: 	jal	yj_fneg
"10101011110111100000000000001111",	-- 8147: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 8148: 	lw	%ra, [%sp + 14]
"10110000000111100000000000001110",	-- 8149: 	sf	%f0, [%sp + 14]
"00111111111111100000000000001111",	-- 8150: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 8151: 	addi	%sp, %sp, 16
"01011000000000000000010011010110",	-- 8152: 	jal	fispos.2522
"10101011110111100000000000010000",	-- 8153: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 8154: 	lw	%ra, [%sp + 15]
"11001100000000100000000000000000",	-- 8155: 	lli	%r2, 0
"00101000001000100000000000000100",	-- 8156: 	bneq	%r1, %r2, bneq_else.9207
"00010100000000000000000000000000",	-- 8157: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 8158: 	lhif	%f0, 0.000000
"01010100000000000001111111100001",	-- 8159: 	j	bneq_cont.9208
	-- bneq_else.9207:
"10010011110000000000000000001110",	-- 8160: 	lf	%f0, [%sp + 14]
	-- bneq_cont.9208:
"10010011110000010000000000000010",	-- 8161: 	lf	%f1, [%sp + 2]
"11101000001000000000000000000000",	-- 8162: 	mulf	%f0, %f1, %f0
"00111011110000010000000000001101",	-- 8163: 	lw	%r1, [%sp + 13]
"10110000000111100000000000001111",	-- 8164: 	sf	%f0, [%sp + 15]
"00111111111111100000000000010000",	-- 8165: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 8166: 	addi	%sp, %sp, 17
"01011000000000000000011001111010",	-- 8167: 	jal	o_diffuse.2646
"10101011110111100000000000010001",	-- 8168: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 8169: 	lw	%ra, [%sp + 16]
"10010011110000010000000000001111",	-- 8170: 	lf	%f1, [%sp + 15]
"11101000001000000000000000000000",	-- 8171: 	mulf	%f0, %f1, %f0
"00111011110000010000000000000001",	-- 8172: 	lw	%r1, [%sp + 1]
"00111011110000100000000000000000",	-- 8173: 	lw	%r2, [%sp + 0]
"01010100000000000000010111001110",	-- 8174: 	j	vecaccum.2605
	-- bneq_else.9206:
"01001111111000000000000000000000",	-- 8175: 	jr	%ra
	-- iter_trace_diffuse_rays.2912:
"00111011011001010000000000000001",	-- 8176: 	lw	%r5, [%r27 + 1]
"11001100000001100000000000000000",	-- 8177: 	lli	%r6, 0
"00110000110001000000000001001000",	-- 8178: 	bgt	%r6, %r4, bgt_else.9210
"10000100001001000011000000000000",	-- 8179: 	add	%r6, %r1, %r4
"00111000110001100000000000000000",	-- 8180: 	lw	%r6, [%r6 + 0]
"00111100011111100000000000000000",	-- 8181: 	sw	%r3, [%sp + 0]
"00111111011111100000000000000001",	-- 8182: 	sw	%r27, [%sp + 1]
"00111100101111100000000000000010",	-- 8183: 	sw	%r5, [%sp + 2]
"00111100100111100000000000000011",	-- 8184: 	sw	%r4, [%sp + 3]
"00111100001111100000000000000100",	-- 8185: 	sw	%r1, [%sp + 4]
"00111100010111100000000000000101",	-- 8186: 	sw	%r2, [%sp + 5]
"10000100000001100000100000000000",	-- 8187: 	add	%r1, %r0, %r6
"00111111111111100000000000000110",	-- 8188: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8189: 	addi	%sp, %sp, 7
"01011000000000000000011010111100",	-- 8190: 	jal	d_vec.2683
"10101011110111100000000000000111",	-- 8191: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8192: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000101",	-- 8193: 	lw	%r2, [%sp + 5]
"00111111111111100000000000000110",	-- 8194: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8195: 	addi	%sp, %sp, 7
"01011000000000000000010110100111",	-- 8196: 	jal	veciprod.2597
"10101011110111100000000000000111",	-- 8197: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8198: 	lw	%ra, [%sp + 6]
"10110000000111100000000000000110",	-- 8199: 	sf	%f0, [%sp + 6]
"00111111111111100000000000000111",	-- 8200: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 8201: 	addi	%sp, %sp, 8
"01011000000000000000010011011101",	-- 8202: 	jal	fisneg.2524
"10101011110111100000000000001000",	-- 8203: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8204: 	lw	%ra, [%sp + 7]
"11001100000000100000000000000000",	-- 8205: 	lli	%r2, 0
"00101000001000100000000000010010",	-- 8206: 	bneq	%r1, %r2, bneq_else.9211
"00111011110000010000000000000011",	-- 8207: 	lw	%r1, [%sp + 3]
"00111011110000100000000000000100",	-- 8208: 	lw	%r2, [%sp + 4]
"10000100010000010001100000000000",	-- 8209: 	add	%r3, %r2, %r1
"00111000011000110000000000000000",	-- 8210: 	lw	%r3, [%r3 + 0]
"00010100000000000000000000000000",	-- 8211: 	llif	%f0, 150.000000
"00010000000000000100001100010110",	-- 8212: 	lhif	%f0, 150.000000
"10010011110000010000000000000110",	-- 8213: 	lf	%f1, [%sp + 6]
"11101100001000000000000000000000",	-- 8214: 	divf	%f0, %f1, %f0
"00111011110110110000000000000010",	-- 8215: 	lw	%r27, [%sp + 2]
"10000100000000110000100000000000",	-- 8216: 	add	%r1, %r0, %r3
"00111111111111100000000000000111",	-- 8217: 	sw	%ra, [%sp + 7]
"00111011011110100000000000000000",	-- 8218: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001000",	-- 8219: 	addi	%sp, %sp, 8
"01010011010000000000000000000000",	-- 8220: 	jalr	%r26
"10101011110111100000000000001000",	-- 8221: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8222: 	lw	%ra, [%sp + 7]
"01010100000000000010000000110001",	-- 8223: 	j	bneq_cont.9212
	-- bneq_else.9211:
"11001100000000010000000000000001",	-- 8224: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 8225: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 8226: 	add	%r1, %r2, %r1
"00111011110000110000000000000100",	-- 8227: 	lw	%r3, [%sp + 4]
"10000100011000010000100000000000",	-- 8228: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 8229: 	lw	%r1, [%r1 + 0]
"00010100000000000000000000000000",	-- 8230: 	llif	%f0, -150.000000
"00010000000000001100001100010110",	-- 8231: 	lhif	%f0, -150.000000
"10010011110000010000000000000110",	-- 8232: 	lf	%f1, [%sp + 6]
"11101100001000000000000000000000",	-- 8233: 	divf	%f0, %f1, %f0
"00111011110110110000000000000010",	-- 8234: 	lw	%r27, [%sp + 2]
"00111111111111100000000000000111",	-- 8235: 	sw	%ra, [%sp + 7]
"00111011011110100000000000000000",	-- 8236: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001000",	-- 8237: 	addi	%sp, %sp, 8
"01010011010000000000000000000000",	-- 8238: 	jalr	%r26
"10101011110111100000000000001000",	-- 8239: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8240: 	lw	%ra, [%sp + 7]
	-- bneq_cont.9212:
"11001100000000010000000000000010",	-- 8241: 	lli	%r1, 2
"00111011110000100000000000000011",	-- 8242: 	lw	%r2, [%sp + 3]
"10001000010000010010000000000000",	-- 8243: 	sub	%r4, %r2, %r1
"00111011110000010000000000000100",	-- 8244: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000101",	-- 8245: 	lw	%r2, [%sp + 5]
"00111011110000110000000000000000",	-- 8246: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000001",	-- 8247: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 8248: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8249: 	jr	%r26
	-- bgt_else.9210:
"01001111111000000000000000000000",	-- 8250: 	jr	%ra
	-- trace_diffuse_rays.2917:
"00111011011001000000000000000010",	-- 8251: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 8252: 	lw	%r5, [%r27 + 1]
"00111100011111100000000000000000",	-- 8253: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 8254: 	sw	%r2, [%sp + 1]
"00111100001111100000000000000010",	-- 8255: 	sw	%r1, [%sp + 2]
"00111100101111100000000000000011",	-- 8256: 	sw	%r5, [%sp + 3]
"10000100000000110000100000000000",	-- 8257: 	add	%r1, %r0, %r3
"10000100000001001101100000000000",	-- 8258: 	add	%r27, %r0, %r4
"00111111111111100000000000000100",	-- 8259: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 8260: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 8261: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 8262: 	jalr	%r26
"10101011110111100000000000000101",	-- 8263: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 8264: 	lw	%ra, [%sp + 4]
"11001100000001000000000001110110",	-- 8265: 	lli	%r4, 118
"00111011110000010000000000000010",	-- 8266: 	lw	%r1, [%sp + 2]
"00111011110000100000000000000001",	-- 8267: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 8268: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000011",	-- 8269: 	lw	%r27, [%sp + 3]
"00111011011110100000000000000000",	-- 8270: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8271: 	jr	%r26
	-- trace_diffuse_ray_80percent.2921:
"00111011011001000000000000000010",	-- 8272: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 8273: 	lw	%r5, [%r27 + 1]
"11001100000001100000000000000000",	-- 8274: 	lli	%r6, 0
"00111100011111100000000000000000",	-- 8275: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 8276: 	sw	%r2, [%sp + 1]
"00111100100111100000000000000010",	-- 8277: 	sw	%r4, [%sp + 2]
"00111100101111100000000000000011",	-- 8278: 	sw	%r5, [%sp + 3]
"00111100001111100000000000000100",	-- 8279: 	sw	%r1, [%sp + 4]
"00101000001001100000000000000010",	-- 8280: 	bneq	%r1, %r6, bneq_else.9214
"01010100000000000010000001100101",	-- 8281: 	j	bneq_cont.9215
	-- bneq_else.9214:
"11001100000001100000000000000000",	-- 8282: 	lli	%r6, 0
"10000100101001100011000000000000",	-- 8283: 	add	%r6, %r5, %r6
"00111000110001100000000000000000",	-- 8284: 	lw	%r6, [%r6 + 0]
"10000100000001100000100000000000",	-- 8285: 	add	%r1, %r0, %r6
"10000100000001001101100000000000",	-- 8286: 	add	%r27, %r0, %r4
"00111111111111100000000000000101",	-- 8287: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 8288: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 8289: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 8290: 	jalr	%r26
"10101011110111100000000000000110",	-- 8291: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 8292: 	lw	%ra, [%sp + 5]
	-- bneq_cont.9215:
"11001100000000010000000000000001",	-- 8293: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 8294: 	lw	%r2, [%sp + 4]
"00101000010000010000000000000010",	-- 8295: 	bneq	%r2, %r1, bneq_else.9216
"01010100000000000010000001111000",	-- 8296: 	j	bneq_cont.9217
	-- bneq_else.9216:
"11001100000000010000000000000001",	-- 8297: 	lli	%r1, 1
"00111011110000110000000000000011",	-- 8298: 	lw	%r3, [%sp + 3]
"10000100011000010000100000000000",	-- 8299: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 8300: 	lw	%r1, [%r1 + 0]
"00111011110001000000000000000001",	-- 8301: 	lw	%r4, [%sp + 1]
"00111011110001010000000000000000",	-- 8302: 	lw	%r5, [%sp + 0]
"00111011110110110000000000000010",	-- 8303: 	lw	%r27, [%sp + 2]
"10000100000001010001100000000000",	-- 8304: 	add	%r3, %r0, %r5
"10000100000001000001000000000000",	-- 8305: 	add	%r2, %r0, %r4
"00111111111111100000000000000101",	-- 8306: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 8307: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 8308: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 8309: 	jalr	%r26
"10101011110111100000000000000110",	-- 8310: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 8311: 	lw	%ra, [%sp + 5]
	-- bneq_cont.9217:
"11001100000000010000000000000010",	-- 8312: 	lli	%r1, 2
"00111011110000100000000000000100",	-- 8313: 	lw	%r2, [%sp + 4]
"00101000010000010000000000000010",	-- 8314: 	bneq	%r2, %r1, bneq_else.9218
"01010100000000000010000010001011",	-- 8315: 	j	bneq_cont.9219
	-- bneq_else.9218:
"11001100000000010000000000000010",	-- 8316: 	lli	%r1, 2
"00111011110000110000000000000011",	-- 8317: 	lw	%r3, [%sp + 3]
"10000100011000010000100000000000",	-- 8318: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 8319: 	lw	%r1, [%r1 + 0]
"00111011110001000000000000000001",	-- 8320: 	lw	%r4, [%sp + 1]
"00111011110001010000000000000000",	-- 8321: 	lw	%r5, [%sp + 0]
"00111011110110110000000000000010",	-- 8322: 	lw	%r27, [%sp + 2]
"10000100000001010001100000000000",	-- 8323: 	add	%r3, %r0, %r5
"10000100000001000001000000000000",	-- 8324: 	add	%r2, %r0, %r4
"00111111111111100000000000000101",	-- 8325: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 8326: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 8327: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 8328: 	jalr	%r26
"10101011110111100000000000000110",	-- 8329: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 8330: 	lw	%ra, [%sp + 5]
	-- bneq_cont.9219:
"11001100000000010000000000000011",	-- 8331: 	lli	%r1, 3
"00111011110000100000000000000100",	-- 8332: 	lw	%r2, [%sp + 4]
"00101000010000010000000000000010",	-- 8333: 	bneq	%r2, %r1, bneq_else.9220
"01010100000000000010000010011110",	-- 8334: 	j	bneq_cont.9221
	-- bneq_else.9220:
"11001100000000010000000000000011",	-- 8335: 	lli	%r1, 3
"00111011110000110000000000000011",	-- 8336: 	lw	%r3, [%sp + 3]
"10000100011000010000100000000000",	-- 8337: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 8338: 	lw	%r1, [%r1 + 0]
"00111011110001000000000000000001",	-- 8339: 	lw	%r4, [%sp + 1]
"00111011110001010000000000000000",	-- 8340: 	lw	%r5, [%sp + 0]
"00111011110110110000000000000010",	-- 8341: 	lw	%r27, [%sp + 2]
"10000100000001010001100000000000",	-- 8342: 	add	%r3, %r0, %r5
"10000100000001000001000000000000",	-- 8343: 	add	%r2, %r0, %r4
"00111111111111100000000000000101",	-- 8344: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 8345: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 8346: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 8347: 	jalr	%r26
"10101011110111100000000000000110",	-- 8348: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 8349: 	lw	%ra, [%sp + 5]
	-- bneq_cont.9221:
"11001100000000010000000000000100",	-- 8350: 	lli	%r1, 4
"00111011110000100000000000000100",	-- 8351: 	lw	%r2, [%sp + 4]
"00101000010000010000000000000010",	-- 8352: 	bneq	%r2, %r1, bneq_else.9222
"01001111111000000000000000000000",	-- 8353: 	jr	%ra
	-- bneq_else.9222:
"11001100000000010000000000000100",	-- 8354: 	lli	%r1, 4
"00111011110000100000000000000011",	-- 8355: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 8356: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8357: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000000001",	-- 8358: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 8359: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000010",	-- 8360: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 8361: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8362: 	jr	%r26
	-- calc_diffuse_using_1point.2925:
"00111011011000110000000000000011",	-- 8363: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 8364: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 8365: 	lw	%r5, [%r27 + 1]
"00111100100111100000000000000000",	-- 8366: 	sw	%r4, [%sp + 0]
"00111100011111100000000000000001",	-- 8367: 	sw	%r3, [%sp + 1]
"00111100101111100000000000000010",	-- 8368: 	sw	%r5, [%sp + 2]
"00111100010111100000000000000011",	-- 8369: 	sw	%r2, [%sp + 3]
"00111100001111100000000000000100",	-- 8370: 	sw	%r1, [%sp + 4]
"00111111111111100000000000000101",	-- 8371: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 8372: 	addi	%sp, %sp, 6
"01011000000000000000011010101110",	-- 8373: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000000110",	-- 8374: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 8375: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000100",	-- 8376: 	lw	%r2, [%sp + 4]
"00111100001111100000000000000101",	-- 8377: 	sw	%r1, [%sp + 5]
"10000100000000100000100000000000",	-- 8378: 	add	%r1, %r0, %r2
"00111111111111100000000000000110",	-- 8379: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8380: 	addi	%sp, %sp, 7
"01011000000000000000011010111010",	-- 8381: 	jal	p_nvectors.2681
"10101011110111100000000000000111",	-- 8382: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8383: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000100",	-- 8384: 	lw	%r2, [%sp + 4]
"00111100001111100000000000000110",	-- 8385: 	sw	%r1, [%sp + 6]
"10000100000000100000100000000000",	-- 8386: 	add	%r1, %r0, %r2
"00111111111111100000000000000111",	-- 8387: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 8388: 	addi	%sp, %sp, 8
"01011000000000000000011010100110",	-- 8389: 	jal	p_intersection_points.2666
"10101011110111100000000000001000",	-- 8390: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8391: 	lw	%ra, [%sp + 7]
"00111011110000100000000000000100",	-- 8392: 	lw	%r2, [%sp + 4]
"00111100001111100000000000000111",	-- 8393: 	sw	%r1, [%sp + 7]
"10000100000000100000100000000000",	-- 8394: 	add	%r1, %r0, %r2
"00111111111111100000000000001000",	-- 8395: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 8396: 	addi	%sp, %sp, 9
"01011000000000000000011010101100",	-- 8397: 	jal	p_energy.2672
"10101011110111100000000000001001",	-- 8398: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 8399: 	lw	%ra, [%sp + 8]
"00111011110000100000000000000011",	-- 8400: 	lw	%r2, [%sp + 3]
"00111011110000110000000000000101",	-- 8401: 	lw	%r3, [%sp + 5]
"10000100011000100001100000000000",	-- 8402: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 8403: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000000010",	-- 8404: 	lw	%r4, [%sp + 2]
"00111100001111100000000000001000",	-- 8405: 	sw	%r1, [%sp + 8]
"10000100000000110001000000000000",	-- 8406: 	add	%r2, %r0, %r3
"10000100000001000000100000000000",	-- 8407: 	add	%r1, %r0, %r4
"00111111111111100000000000001001",	-- 8408: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 8409: 	addi	%sp, %sp, 10
"01011000000000000000010100111101",	-- 8410: 	jal	veccpy.2586
"10101011110111100000000000001010",	-- 8411: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 8412: 	lw	%ra, [%sp + 9]
"00111011110000010000000000000100",	-- 8413: 	lw	%r1, [%sp + 4]
"00111111111111100000000000001001",	-- 8414: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 8415: 	addi	%sp, %sp, 10
"01011000000000000000011010110000",	-- 8416: 	jal	p_group_id.2676
"10101011110111100000000000001010",	-- 8417: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 8418: 	lw	%ra, [%sp + 9]
"00111011110000100000000000000011",	-- 8419: 	lw	%r2, [%sp + 3]
"00111011110000110000000000000110",	-- 8420: 	lw	%r3, [%sp + 6]
"10000100011000100001100000000000",	-- 8421: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 8422: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000000111",	-- 8423: 	lw	%r4, [%sp + 7]
"10000100100000100010000000000000",	-- 8424: 	add	%r4, %r4, %r2
"00111000100001000000000000000000",	-- 8425: 	lw	%r4, [%r4 + 0]
"00111011110110110000000000000001",	-- 8426: 	lw	%r27, [%sp + 1]
"10000100000000110001000000000000",	-- 8427: 	add	%r2, %r0, %r3
"10000100000001000001100000000000",	-- 8428: 	add	%r3, %r0, %r4
"00111111111111100000000000001001",	-- 8429: 	sw	%ra, [%sp + 9]
"00111011011110100000000000000000",	-- 8430: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001010",	-- 8431: 	addi	%sp, %sp, 10
"01010011010000000000000000000000",	-- 8432: 	jalr	%r26
"10101011110111100000000000001010",	-- 8433: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 8434: 	lw	%ra, [%sp + 9]
"00111011110000010000000000000011",	-- 8435: 	lw	%r1, [%sp + 3]
"00111011110000100000000000001000",	-- 8436: 	lw	%r2, [%sp + 8]
"10000100010000010000100000000000",	-- 8437: 	add	%r1, %r2, %r1
"00111000001000100000000000000000",	-- 8438: 	lw	%r2, [%r1 + 0]
"00111011110000010000000000000000",	-- 8439: 	lw	%r1, [%sp + 0]
"00111011110000110000000000000010",	-- 8440: 	lw	%r3, [%sp + 2]
"01010100000000000000011000100101",	-- 8441: 	j	vecaccumv.2618
	-- calc_diffuse_using_5points.2928:
"00111011011001100000000000000010",	-- 8442: 	lw	%r6, [%r27 + 2]
"00111011011001110000000000000001",	-- 8443: 	lw	%r7, [%r27 + 1]
"10000100010000010001000000000000",	-- 8444: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 8445: 	lw	%r2, [%r2 + 0]
"00111100110111100000000000000000",	-- 8446: 	sw	%r6, [%sp + 0]
"00111100111111100000000000000001",	-- 8447: 	sw	%r7, [%sp + 1]
"00111100101111100000000000000010",	-- 8448: 	sw	%r5, [%sp + 2]
"00111100100111100000000000000011",	-- 8449: 	sw	%r4, [%sp + 3]
"00111100011111100000000000000100",	-- 8450: 	sw	%r3, [%sp + 4]
"00111100001111100000000000000101",	-- 8451: 	sw	%r1, [%sp + 5]
"10000100000000100000100000000000",	-- 8452: 	add	%r1, %r0, %r2
"00111111111111100000000000000110",	-- 8453: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8454: 	addi	%sp, %sp, 7
"01011000000000000000011010101110",	-- 8455: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000000111",	-- 8456: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8457: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000001",	-- 8458: 	lli	%r2, 1
"00111011110000110000000000000101",	-- 8459: 	lw	%r3, [%sp + 5]
"10001000011000100001000000000000",	-- 8460: 	sub	%r2, %r3, %r2
"00111011110001000000000000000100",	-- 8461: 	lw	%r4, [%sp + 4]
"10000100100000100001000000000000",	-- 8462: 	add	%r2, %r4, %r2
"00111000010000100000000000000000",	-- 8463: 	lw	%r2, [%r2 + 0]
"00111100001111100000000000000110",	-- 8464: 	sw	%r1, [%sp + 6]
"10000100000000100000100000000000",	-- 8465: 	add	%r1, %r0, %r2
"00111111111111100000000000000111",	-- 8466: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 8467: 	addi	%sp, %sp, 8
"01011000000000000000011010101110",	-- 8468: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000001000",	-- 8469: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8470: 	lw	%ra, [%sp + 7]
"00111011110000100000000000000101",	-- 8471: 	lw	%r2, [%sp + 5]
"00111011110000110000000000000100",	-- 8472: 	lw	%r3, [%sp + 4]
"10000100011000100010000000000000",	-- 8473: 	add	%r4, %r3, %r2
"00111000100001000000000000000000",	-- 8474: 	lw	%r4, [%r4 + 0]
"00111100001111100000000000000111",	-- 8475: 	sw	%r1, [%sp + 7]
"10000100000001000000100000000000",	-- 8476: 	add	%r1, %r0, %r4
"00111111111111100000000000001000",	-- 8477: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 8478: 	addi	%sp, %sp, 9
"01011000000000000000011010101110",	-- 8479: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000001001",	-- 8480: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 8481: 	lw	%ra, [%sp + 8]
"11001100000000100000000000000001",	-- 8482: 	lli	%r2, 1
"00111011110000110000000000000101",	-- 8483: 	lw	%r3, [%sp + 5]
"10000100011000100001000000000000",	-- 8484: 	add	%r2, %r3, %r2
"00111011110001000000000000000100",	-- 8485: 	lw	%r4, [%sp + 4]
"10000100100000100001000000000000",	-- 8486: 	add	%r2, %r4, %r2
"00111000010000100000000000000000",	-- 8487: 	lw	%r2, [%r2 + 0]
"00111100001111100000000000001000",	-- 8488: 	sw	%r1, [%sp + 8]
"10000100000000100000100000000000",	-- 8489: 	add	%r1, %r0, %r2
"00111111111111100000000000001001",	-- 8490: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 8491: 	addi	%sp, %sp, 10
"01011000000000000000011010101110",	-- 8492: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000001010",	-- 8493: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 8494: 	lw	%ra, [%sp + 9]
"00111011110000100000000000000101",	-- 8495: 	lw	%r2, [%sp + 5]
"00111011110000110000000000000011",	-- 8496: 	lw	%r3, [%sp + 3]
"10000100011000100001100000000000",	-- 8497: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 8498: 	lw	%r3, [%r3 + 0]
"00111100001111100000000000001001",	-- 8499: 	sw	%r1, [%sp + 9]
"10000100000000110000100000000000",	-- 8500: 	add	%r1, %r0, %r3
"00111111111111100000000000001010",	-- 8501: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 8502: 	addi	%sp, %sp, 11
"01011000000000000000011010101110",	-- 8503: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000001011",	-- 8504: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 8505: 	lw	%ra, [%sp + 10]
"00111011110000100000000000000010",	-- 8506: 	lw	%r2, [%sp + 2]
"00111011110000110000000000000110",	-- 8507: 	lw	%r3, [%sp + 6]
"10000100011000100001100000000000",	-- 8508: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 8509: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000000001",	-- 8510: 	lw	%r4, [%sp + 1]
"00111100001111100000000000001010",	-- 8511: 	sw	%r1, [%sp + 10]
"10000100000000110001000000000000",	-- 8512: 	add	%r2, %r0, %r3
"10000100000001000000100000000000",	-- 8513: 	add	%r1, %r0, %r4
"00111111111111100000000000001011",	-- 8514: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8515: 	addi	%sp, %sp, 12
"01011000000000000000010100111101",	-- 8516: 	jal	veccpy.2586
"10101011110111100000000000001100",	-- 8517: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8518: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000010",	-- 8519: 	lw	%r1, [%sp + 2]
"00111011110000100000000000000111",	-- 8520: 	lw	%r2, [%sp + 7]
"10000100010000010001000000000000",	-- 8521: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 8522: 	lw	%r2, [%r2 + 0]
"00111011110000110000000000000001",	-- 8523: 	lw	%r3, [%sp + 1]
"10000100000000110000100000000000",	-- 8524: 	add	%r1, %r0, %r3
"00111111111111100000000000001011",	-- 8525: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8526: 	addi	%sp, %sp, 12
"01011000000000000000010111110000",	-- 8527: 	jal	vecadd.2609
"10101011110111100000000000001100",	-- 8528: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8529: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000010",	-- 8530: 	lw	%r1, [%sp + 2]
"00111011110000100000000000001000",	-- 8531: 	lw	%r2, [%sp + 8]
"10000100010000010001000000000000",	-- 8532: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 8533: 	lw	%r2, [%r2 + 0]
"00111011110000110000000000000001",	-- 8534: 	lw	%r3, [%sp + 1]
"10000100000000110000100000000000",	-- 8535: 	add	%r1, %r0, %r3
"00111111111111100000000000001011",	-- 8536: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8537: 	addi	%sp, %sp, 12
"01011000000000000000010111110000",	-- 8538: 	jal	vecadd.2609
"10101011110111100000000000001100",	-- 8539: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8540: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000010",	-- 8541: 	lw	%r1, [%sp + 2]
"00111011110000100000000000001001",	-- 8542: 	lw	%r2, [%sp + 9]
"10000100010000010001000000000000",	-- 8543: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 8544: 	lw	%r2, [%r2 + 0]
"00111011110000110000000000000001",	-- 8545: 	lw	%r3, [%sp + 1]
"10000100000000110000100000000000",	-- 8546: 	add	%r1, %r0, %r3
"00111111111111100000000000001011",	-- 8547: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8548: 	addi	%sp, %sp, 12
"01011000000000000000010111110000",	-- 8549: 	jal	vecadd.2609
"10101011110111100000000000001100",	-- 8550: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8551: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000010",	-- 8552: 	lw	%r1, [%sp + 2]
"00111011110000100000000000001010",	-- 8553: 	lw	%r2, [%sp + 10]
"10000100010000010001000000000000",	-- 8554: 	add	%r2, %r2, %r1
"00111000010000100000000000000000",	-- 8555: 	lw	%r2, [%r2 + 0]
"00111011110000110000000000000001",	-- 8556: 	lw	%r3, [%sp + 1]
"10000100000000110000100000000000",	-- 8557: 	add	%r1, %r0, %r3
"00111111111111100000000000001011",	-- 8558: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8559: 	addi	%sp, %sp, 12
"01011000000000000000010111110000",	-- 8560: 	jal	vecadd.2609
"10101011110111100000000000001100",	-- 8561: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8562: 	lw	%ra, [%sp + 11]
"00111011110000010000000000000101",	-- 8563: 	lw	%r1, [%sp + 5]
"00111011110000100000000000000100",	-- 8564: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 8565: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8566: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001011",	-- 8567: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8568: 	addi	%sp, %sp, 12
"01011000000000000000011010101100",	-- 8569: 	jal	p_energy.2672
"10101011110111100000000000001100",	-- 8570: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8571: 	lw	%ra, [%sp + 11]
"00111011110000100000000000000010",	-- 8572: 	lw	%r2, [%sp + 2]
"10000100001000100000100000000000",	-- 8573: 	add	%r1, %r1, %r2
"00111000001000100000000000000000",	-- 8574: 	lw	%r2, [%r1 + 0]
"00111011110000010000000000000000",	-- 8575: 	lw	%r1, [%sp + 0]
"00111011110000110000000000000001",	-- 8576: 	lw	%r3, [%sp + 1]
"01010100000000000000011000100101",	-- 8577: 	j	vecaccumv.2618
	-- do_without_neighbors.2934:
"00111011011000110000000000000001",	-- 8578: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000100",	-- 8579: 	lli	%r4, 4
"00110000010001000000000000101011",	-- 8580: 	bgt	%r2, %r4, bgt_else.9224
"00111111011111100000000000000000",	-- 8581: 	sw	%r27, [%sp + 0]
"00111100011111100000000000000001",	-- 8582: 	sw	%r3, [%sp + 1]
"00111100001111100000000000000010",	-- 8583: 	sw	%r1, [%sp + 2]
"00111100010111100000000000000011",	-- 8584: 	sw	%r2, [%sp + 3]
"00111111111111100000000000000100",	-- 8585: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 8586: 	addi	%sp, %sp, 5
"01011000000000000000011010101000",	-- 8587: 	jal	p_surface_ids.2668
"10101011110111100000000000000101",	-- 8588: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 8589: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000000",	-- 8590: 	lli	%r2, 0
"00111011110000110000000000000011",	-- 8591: 	lw	%r3, [%sp + 3]
"10000100001000110000100000000000",	-- 8592: 	add	%r1, %r1, %r3
"00111000001000010000000000000000",	-- 8593: 	lw	%r1, [%r1 + 0]
"00110000010000010000000000011100",	-- 8594: 	bgt	%r2, %r1, bgt_else.9225
"00111011110000010000000000000010",	-- 8595: 	lw	%r1, [%sp + 2]
"00111111111111100000000000000100",	-- 8596: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 8597: 	addi	%sp, %sp, 5
"01011000000000000000011010101010",	-- 8598: 	jal	p_calc_diffuse.2670
"10101011110111100000000000000101",	-- 8599: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 8600: 	lw	%ra, [%sp + 4]
"00111011110000100000000000000011",	-- 8601: 	lw	%r2, [%sp + 3]
"10000100001000100000100000000000",	-- 8602: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 8603: 	lw	%r1, [%r1 + 0]
"11001100000000110000000000000000",	-- 8604: 	lli	%r3, 0
"00101000001000110000000000000010",	-- 8605: 	bneq	%r1, %r3, bneq_else.9226
"01010100000000000010000110100111",	-- 8606: 	j	bneq_cont.9227
	-- bneq_else.9226:
"00111011110000010000000000000010",	-- 8607: 	lw	%r1, [%sp + 2]
"00111011110110110000000000000001",	-- 8608: 	lw	%r27, [%sp + 1]
"00111111111111100000000000000100",	-- 8609: 	sw	%ra, [%sp + 4]
"00111011011110100000000000000000",	-- 8610: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000101",	-- 8611: 	addi	%sp, %sp, 5
"01010011010000000000000000000000",	-- 8612: 	jalr	%r26
"10101011110111100000000000000101",	-- 8613: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 8614: 	lw	%ra, [%sp + 4]
	-- bneq_cont.9227:
"11001100000000010000000000000001",	-- 8615: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 8616: 	lw	%r2, [%sp + 3]
"10000100010000010001000000000000",	-- 8617: 	add	%r2, %r2, %r1
"00111011110000010000000000000010",	-- 8618: 	lw	%r1, [%sp + 2]
"00111011110110110000000000000000",	-- 8619: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 8620: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8621: 	jr	%r26
	-- bgt_else.9225:
"01001111111000000000000000000000",	-- 8622: 	jr	%ra
	-- bgt_else.9224:
"01001111111000000000000000000000",	-- 8623: 	jr	%ra
	-- neighbors_exist.2937:
"00111011011000110000000000000001",	-- 8624: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000001",	-- 8625: 	lli	%r4, 1
"10000100011001000010000000000000",	-- 8626: 	add	%r4, %r3, %r4
"00111000100001000000000000000000",	-- 8627: 	lw	%r4, [%r4 + 0]
"11001100000001010000000000000001",	-- 8628: 	lli	%r5, 1
"10000100010001010010100000000000",	-- 8629: 	add	%r5, %r2, %r5
"00110000100001010000000000000011",	-- 8630: 	bgt	%r4, %r5, bgt_else.9230
"11001100000000010000000000000000",	-- 8631: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8632: 	jr	%ra
	-- bgt_else.9230:
"11001100000001000000000000000000",	-- 8633: 	lli	%r4, 0
"00110000010001000000000000000011",	-- 8634: 	bgt	%r2, %r4, bgt_else.9231
"11001100000000010000000000000000",	-- 8635: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8636: 	jr	%ra
	-- bgt_else.9231:
"11001100000000100000000000000000",	-- 8637: 	lli	%r2, 0
"10000100011000100001000000000000",	-- 8638: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 8639: 	lw	%r2, [%r2 + 0]
"11001100000000110000000000000001",	-- 8640: 	lli	%r3, 1
"10000100001000110001100000000000",	-- 8641: 	add	%r3, %r1, %r3
"00110000010000110000000000000011",	-- 8642: 	bgt	%r2, %r3, bgt_else.9232
"11001100000000010000000000000000",	-- 8643: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8644: 	jr	%ra
	-- bgt_else.9232:
"11001100000000100000000000000000",	-- 8645: 	lli	%r2, 0
"00110000001000100000000000000011",	-- 8646: 	bgt	%r1, %r2, bgt_else.9233
"11001100000000010000000000000000",	-- 8647: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8648: 	jr	%ra
	-- bgt_else.9233:
"11001100000000010000000000000001",	-- 8649: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 8650: 	jr	%ra
	-- get_surface_id.2941:
"00111100010111100000000000000000",	-- 8651: 	sw	%r2, [%sp + 0]
"00111111111111100000000000000001",	-- 8652: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8653: 	addi	%sp, %sp, 2
"01011000000000000000011010101000",	-- 8654: 	jal	p_surface_ids.2668
"10101011110111100000000000000010",	-- 8655: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8656: 	lw	%ra, [%sp + 1]
"00111011110000100000000000000000",	-- 8657: 	lw	%r2, [%sp + 0]
"10000100001000100000100000000000",	-- 8658: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 8659: 	lw	%r1, [%r1 + 0]
"01001111111000000000000000000000",	-- 8660: 	jr	%ra
	-- neighbors_are_available.2944:
"10000100011000010011000000000000",	-- 8661: 	add	%r6, %r3, %r1
"00111000110001100000000000000000",	-- 8662: 	lw	%r6, [%r6 + 0]
"00111100011111100000000000000000",	-- 8663: 	sw	%r3, [%sp + 0]
"00111100100111100000000000000001",	-- 8664: 	sw	%r4, [%sp + 1]
"00111100101111100000000000000010",	-- 8665: 	sw	%r5, [%sp + 2]
"00111100001111100000000000000011",	-- 8666: 	sw	%r1, [%sp + 3]
"00111100010111100000000000000100",	-- 8667: 	sw	%r2, [%sp + 4]
"10000100000001010001000000000000",	-- 8668: 	add	%r2, %r0, %r5
"10000100000001100000100000000000",	-- 8669: 	add	%r1, %r0, %r6
"00111111111111100000000000000101",	-- 8670: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 8671: 	addi	%sp, %sp, 6
"01011000000000000010000111001011",	-- 8672: 	jal	get_surface_id.2941
"10101011110111100000000000000110",	-- 8673: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 8674: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000011",	-- 8675: 	lw	%r2, [%sp + 3]
"00111011110000110000000000000100",	-- 8676: 	lw	%r3, [%sp + 4]
"10000100011000100001100000000000",	-- 8677: 	add	%r3, %r3, %r2
"00111000011000110000000000000000",	-- 8678: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000000010",	-- 8679: 	lw	%r4, [%sp + 2]
"00111100001111100000000000000101",	-- 8680: 	sw	%r1, [%sp + 5]
"10000100000001000001000000000000",	-- 8681: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 8682: 	add	%r1, %r0, %r3
"00111111111111100000000000000110",	-- 8683: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8684: 	addi	%sp, %sp, 7
"01011000000000000010000111001011",	-- 8685: 	jal	get_surface_id.2941
"10101011110111100000000000000111",	-- 8686: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8687: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000101",	-- 8688: 	lw	%r2, [%sp + 5]
"00101000001000100000000000110101",	-- 8689: 	bneq	%r1, %r2, bneq_else.9234
"00111011110000010000000000000011",	-- 8690: 	lw	%r1, [%sp + 3]
"00111011110000110000000000000001",	-- 8691: 	lw	%r3, [%sp + 1]
"10000100011000010001100000000000",	-- 8692: 	add	%r3, %r3, %r1
"00111000011000110000000000000000",	-- 8693: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000000010",	-- 8694: 	lw	%r4, [%sp + 2]
"10000100000001000001000000000000",	-- 8695: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 8696: 	add	%r1, %r0, %r3
"00111111111111100000000000000110",	-- 8697: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8698: 	addi	%sp, %sp, 7
"01011000000000000010000111001011",	-- 8699: 	jal	get_surface_id.2941
"10101011110111100000000000000111",	-- 8700: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8701: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000101",	-- 8702: 	lw	%r2, [%sp + 5]
"00101000001000100000000000100101",	-- 8703: 	bneq	%r1, %r2, bneq_else.9235
"11001100000000010000000000000001",	-- 8704: 	lli	%r1, 1
"00111011110000110000000000000011",	-- 8705: 	lw	%r3, [%sp + 3]
"10001000011000010000100000000000",	-- 8706: 	sub	%r1, %r3, %r1
"00111011110001000000000000000000",	-- 8707: 	lw	%r4, [%sp + 0]
"10000100100000010000100000000000",	-- 8708: 	add	%r1, %r4, %r1
"00111000001000010000000000000000",	-- 8709: 	lw	%r1, [%r1 + 0]
"00111011110001010000000000000010",	-- 8710: 	lw	%r5, [%sp + 2]
"10000100000001010001000000000000",	-- 8711: 	add	%r2, %r0, %r5
"00111111111111100000000000000110",	-- 8712: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8713: 	addi	%sp, %sp, 7
"01011000000000000010000111001011",	-- 8714: 	jal	get_surface_id.2941
"10101011110111100000000000000111",	-- 8715: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8716: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000101",	-- 8717: 	lw	%r2, [%sp + 5]
"00101000001000100000000000010100",	-- 8718: 	bneq	%r1, %r2, bneq_else.9236
"11001100000000010000000000000001",	-- 8719: 	lli	%r1, 1
"00111011110000110000000000000011",	-- 8720: 	lw	%r3, [%sp + 3]
"10000100011000010000100000000000",	-- 8721: 	add	%r1, %r3, %r1
"00111011110000110000000000000000",	-- 8722: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 8723: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 8724: 	lw	%r1, [%r1 + 0]
"00111011110000110000000000000010",	-- 8725: 	lw	%r3, [%sp + 2]
"10000100000000110001000000000000",	-- 8726: 	add	%r2, %r0, %r3
"00111111111111100000000000000110",	-- 8727: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8728: 	addi	%sp, %sp, 7
"01011000000000000010000111001011",	-- 8729: 	jal	get_surface_id.2941
"10101011110111100000000000000111",	-- 8730: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8731: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000101",	-- 8732: 	lw	%r2, [%sp + 5]
"00101000001000100000000000000011",	-- 8733: 	bneq	%r1, %r2, bneq_else.9237
"11001100000000010000000000000001",	-- 8734: 	lli	%r1, 1
"01001111111000000000000000000000",	-- 8735: 	jr	%ra
	-- bneq_else.9237:
"11001100000000010000000000000000",	-- 8736: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8737: 	jr	%ra
	-- bneq_else.9236:
"11001100000000010000000000000000",	-- 8738: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8739: 	jr	%ra
	-- bneq_else.9235:
"11001100000000010000000000000000",	-- 8740: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8741: 	jr	%ra
	-- bneq_else.9234:
"11001100000000010000000000000000",	-- 8742: 	lli	%r1, 0
"01001111111000000000000000000000",	-- 8743: 	jr	%ra
	-- try_exploit_neighbors.2950:
"00111011011001110000000000000010",	-- 8744: 	lw	%r7, [%r27 + 2]
"00111011011010000000000000000001",	-- 8745: 	lw	%r8, [%r27 + 1]
"10000100100000010100100000000000",	-- 8746: 	add	%r9, %r4, %r1
"00111001001010010000000000000000",	-- 8747: 	lw	%r9, [%r9 + 0]
"11001100000010100000000000000100",	-- 8748: 	lli	%r10, 4
"00110000110010100000000001001101",	-- 8749: 	bgt	%r6, %r10, bgt_else.9238
"11001100000010100000000000000000",	-- 8750: 	lli	%r10, 0
"00111100010111100000000000000000",	-- 8751: 	sw	%r2, [%sp + 0]
"00111111011111100000000000000001",	-- 8752: 	sw	%r27, [%sp + 1]
"00111101000111100000000000000010",	-- 8753: 	sw	%r8, [%sp + 2]
"00111101001111100000000000000011",	-- 8754: 	sw	%r9, [%sp + 3]
"00111100111111100000000000000100",	-- 8755: 	sw	%r7, [%sp + 4]
"00111100110111100000000000000101",	-- 8756: 	sw	%r6, [%sp + 5]
"00111100101111100000000000000110",	-- 8757: 	sw	%r5, [%sp + 6]
"00111100100111100000000000000111",	-- 8758: 	sw	%r4, [%sp + 7]
"00111100011111100000000000001000",	-- 8759: 	sw	%r3, [%sp + 8]
"00111100001111100000000000001001",	-- 8760: 	sw	%r1, [%sp + 9]
"00111101010111100000000000001010",	-- 8761: 	sw	%r10, [%sp + 10]
"10000100000001100001000000000000",	-- 8762: 	add	%r2, %r0, %r6
"10000100000010010000100000000000",	-- 8763: 	add	%r1, %r0, %r9
"00111111111111100000000000001011",	-- 8764: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8765: 	addi	%sp, %sp, 12
"01011000000000000010000111001011",	-- 8766: 	jal	get_surface_id.2941
"10101011110111100000000000001100",	-- 8767: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8768: 	lw	%ra, [%sp + 11]
"00111011110000100000000000001010",	-- 8769: 	lw	%r2, [%sp + 10]
"00110000010000010000000000110111",	-- 8770: 	bgt	%r2, %r1, bgt_else.9239
"00111011110000010000000000001001",	-- 8771: 	lw	%r1, [%sp + 9]
"00111011110000100000000000001000",	-- 8772: 	lw	%r2, [%sp + 8]
"00111011110000110000000000000111",	-- 8773: 	lw	%r3, [%sp + 7]
"00111011110001000000000000000110",	-- 8774: 	lw	%r4, [%sp + 6]
"00111011110001010000000000000101",	-- 8775: 	lw	%r5, [%sp + 5]
"00111111111111100000000000001011",	-- 8776: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8777: 	addi	%sp, %sp, 12
"01011000000000000010000111010101",	-- 8778: 	jal	neighbors_are_available.2944
"10101011110111100000000000001100",	-- 8779: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8780: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 8781: 	lli	%r2, 0
"00101000001000100000000000001001",	-- 8782: 	bneq	%r1, %r2, bneq_else.9240
"00111011110000010000000000001001",	-- 8783: 	lw	%r1, [%sp + 9]
"00111011110000100000000000000111",	-- 8784: 	lw	%r2, [%sp + 7]
"10000100010000010000100000000000",	-- 8785: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8786: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000000101",	-- 8787: 	lw	%r2, [%sp + 5]
"00111011110110110000000000000100",	-- 8788: 	lw	%r27, [%sp + 4]
"00111011011110100000000000000000",	-- 8789: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8790: 	jr	%r26
	-- bneq_else.9240:
"00111011110000010000000000000011",	-- 8791: 	lw	%r1, [%sp + 3]
"00111111111111100000000000001011",	-- 8792: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 8793: 	addi	%sp, %sp, 12
"01011000000000000000011010101010",	-- 8794: 	jal	p_calc_diffuse.2670
"10101011110111100000000000001100",	-- 8795: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8796: 	lw	%ra, [%sp + 11]
"00111011110001010000000000000101",	-- 8797: 	lw	%r5, [%sp + 5]
"10000100001001010000100000000000",	-- 8798: 	add	%r1, %r1, %r5
"00111000001000010000000000000000",	-- 8799: 	lw	%r1, [%r1 + 0]
"11001100000000100000000000000000",	-- 8800: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 8801: 	bneq	%r1, %r2, bneq_else.9241
"01010100000000000010001001101110",	-- 8802: 	j	bneq_cont.9242
	-- bneq_else.9241:
"00111011110000010000000000001001",	-- 8803: 	lw	%r1, [%sp + 9]
"00111011110000100000000000001000",	-- 8804: 	lw	%r2, [%sp + 8]
"00111011110000110000000000000111",	-- 8805: 	lw	%r3, [%sp + 7]
"00111011110001000000000000000110",	-- 8806: 	lw	%r4, [%sp + 6]
"00111011110110110000000000000010",	-- 8807: 	lw	%r27, [%sp + 2]
"00111111111111100000000000001011",	-- 8808: 	sw	%ra, [%sp + 11]
"00111011011110100000000000000000",	-- 8809: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001100",	-- 8810: 	addi	%sp, %sp, 12
"01010011010000000000000000000000",	-- 8811: 	jalr	%r26
"10101011110111100000000000001100",	-- 8812: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 8813: 	lw	%ra, [%sp + 11]
	-- bneq_cont.9242:
"11001100000000010000000000000001",	-- 8814: 	lli	%r1, 1
"00111011110000100000000000000101",	-- 8815: 	lw	%r2, [%sp + 5]
"10000100010000010011000000000000",	-- 8816: 	add	%r6, %r2, %r1
"00111011110000010000000000001001",	-- 8817: 	lw	%r1, [%sp + 9]
"00111011110000100000000000000000",	-- 8818: 	lw	%r2, [%sp + 0]
"00111011110000110000000000001000",	-- 8819: 	lw	%r3, [%sp + 8]
"00111011110001000000000000000111",	-- 8820: 	lw	%r4, [%sp + 7]
"00111011110001010000000000000110",	-- 8821: 	lw	%r5, [%sp + 6]
"00111011110110110000000000000001",	-- 8822: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 8823: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 8824: 	jr	%r26
	-- bgt_else.9239:
"01001111111000000000000000000000",	-- 8825: 	jr	%ra
	-- bgt_else.9238:
"01001111111000000000000000000000",	-- 8826: 	jr	%ra
	-- write_ppm_header.2957:
"00111011011000010000000000000001",	-- 8827: 	lw	%r1, [%r27 + 1]
"11001100000000100000000001010000",	-- 8828: 	lli	%r2, 80
"00111100001111100000000000000000",	-- 8829: 	sw	%r1, [%sp + 0]
"10000100000000100000100000000000",	-- 8830: 	add	%r1, %r0, %r2
"00111111111111100000000000000001",	-- 8831: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8832: 	addi	%sp, %sp, 2
"01011000000000000010101000011010",	-- 8833: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8834: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8835: 	lw	%ra, [%sp + 1]
"11001100000000010000000000110011",	-- 8836: 	lli	%r1, 51
"00111111111111100000000000000001",	-- 8837: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8838: 	addi	%sp, %sp, 2
"01011000000000000010101000011010",	-- 8839: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8840: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8841: 	lw	%ra, [%sp + 1]
"11001100000000010000000000001010",	-- 8842: 	lli	%r1, 10
"00111111111111100000000000000001",	-- 8843: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8844: 	addi	%sp, %sp, 2
"01011000000000000010101000011010",	-- 8845: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8846: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8847: 	lw	%ra, [%sp + 1]
"11001100000000010000000000000000",	-- 8848: 	lli	%r1, 0
"00111011110000100000000000000000",	-- 8849: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 8850: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8851: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000000001",	-- 8852: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8853: 	addi	%sp, %sp, 2
"01011000000000000000010000000010",	-- 8854: 	jal	print_int.2514
"10101011110111100000000000000010",	-- 8855: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8856: 	lw	%ra, [%sp + 1]
"11001100000000010000000000100000",	-- 8857: 	lli	%r1, 32
"00111111111111100000000000000001",	-- 8858: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8859: 	addi	%sp, %sp, 2
"01011000000000000010101000011010",	-- 8860: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8861: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8862: 	lw	%ra, [%sp + 1]
"11001100000000010000000000000001",	-- 8863: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 8864: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 8865: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 8866: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000000001",	-- 8867: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8868: 	addi	%sp, %sp, 2
"01011000000000000000010000000010",	-- 8869: 	jal	print_int.2514
"10101011110111100000000000000010",	-- 8870: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8871: 	lw	%ra, [%sp + 1]
"11001100000000010000000000100000",	-- 8872: 	lli	%r1, 32
"00111111111111100000000000000001",	-- 8873: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8874: 	addi	%sp, %sp, 2
"01011000000000000010101000011010",	-- 8875: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8876: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8877: 	lw	%ra, [%sp + 1]
"11001100000000010000000011111111",	-- 8878: 	lli	%r1, 255
"00111111111111100000000000000001",	-- 8879: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8880: 	addi	%sp, %sp, 2
"01011000000000000000010000000010",	-- 8881: 	jal	print_int.2514
"10101011110111100000000000000010",	-- 8882: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8883: 	lw	%ra, [%sp + 1]
"11001100000000010000000000001010",	-- 8884: 	lli	%r1, 10
"01010100000000000010101000011010",	-- 8885: 	j	yj_print_char
	-- write_rgb_element.2959:
"00111111111111100000000000000000",	-- 8886: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 8887: 	addi	%sp, %sp, 1
"01011000000000000010101000101110",	-- 8888: 	jal	yj_int_of_float
"10101011110111100000000000000001",	-- 8889: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 8890: 	lw	%ra, [%sp + 0]
"11001100000000100000000011111111",	-- 8891: 	lli	%r2, 255
"00110000001000100000000000000110",	-- 8892: 	bgt	%r1, %r2, bgt_else.9245
"11001100000000100000000000000000",	-- 8893: 	lli	%r2, 0
"00110000010000010000000000000010",	-- 8894: 	bgt	%r2, %r1, bgt_else.9247
"01010100000000000010001011000001",	-- 8895: 	j	bgt_cont.9248
	-- bgt_else.9247:
"11001100000000010000000000000000",	-- 8896: 	lli	%r1, 0
	-- bgt_cont.9248:
"01010100000000000010001011000011",	-- 8897: 	j	bgt_cont.9246
	-- bgt_else.9245:
"11001100000000010000000011111111",	-- 8898: 	lli	%r1, 255
	-- bgt_cont.9246:
"01010100000000000000010000000010",	-- 8899: 	j	print_int.2514
	-- write_rgb.2961:
"00111011011000010000000000000001",	-- 8900: 	lw	%r1, [%r27 + 1]
"11001100000000100000000000000000",	-- 8901: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 8902: 	add	%r2, %r1, %r2
"10010000010000000000000000000000",	-- 8903: 	lf	%f0, [%r2 + 0]
"00111100001111100000000000000000",	-- 8904: 	sw	%r1, [%sp + 0]
"00111111111111100000000000000001",	-- 8905: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8906: 	addi	%sp, %sp, 2
"01011000000000000010001010110110",	-- 8907: 	jal	write_rgb_element.2959
"10101011110111100000000000000010",	-- 8908: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8909: 	lw	%ra, [%sp + 1]
"11001100000000010000000000100000",	-- 8910: 	lli	%r1, 32
"00111111111111100000000000000001",	-- 8911: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8912: 	addi	%sp, %sp, 2
"01011000000000000010101000011010",	-- 8913: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8914: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8915: 	lw	%ra, [%sp + 1]
"11001100000000010000000000000001",	-- 8916: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 8917: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 8918: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 8919: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000000001",	-- 8920: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8921: 	addi	%sp, %sp, 2
"01011000000000000010001010110110",	-- 8922: 	jal	write_rgb_element.2959
"10101011110111100000000000000010",	-- 8923: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8924: 	lw	%ra, [%sp + 1]
"11001100000000010000000000100000",	-- 8925: 	lli	%r1, 32
"00111111111111100000000000000001",	-- 8926: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8927: 	addi	%sp, %sp, 2
"01011000000000000010101000011010",	-- 8928: 	jal	yj_print_char
"10101011110111100000000000000010",	-- 8929: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8930: 	lw	%ra, [%sp + 1]
"11001100000000010000000000000010",	-- 8931: 	lli	%r1, 2
"00111011110000100000000000000000",	-- 8932: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 8933: 	add	%r1, %r2, %r1
"10010000001000000000000000000000",	-- 8934: 	lf	%f0, [%r1 + 0]
"00111111111111100000000000000001",	-- 8935: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 8936: 	addi	%sp, %sp, 2
"01011000000000000010001010110110",	-- 8937: 	jal	write_rgb_element.2959
"10101011110111100000000000000010",	-- 8938: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 8939: 	lw	%ra, [%sp + 1]
"11001100000000010000000000001010",	-- 8940: 	lli	%r1, 10
"01010100000000000010101000011010",	-- 8941: 	j	yj_print_char
	-- pretrace_diffuse_rays.2963:
"00111011011000110000000000000011",	-- 8942: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 8943: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 8944: 	lw	%r5, [%r27 + 1]
"11001100000001100000000000000100",	-- 8945: 	lli	%r6, 4
"00110000010001100000000001100010",	-- 8946: 	bgt	%r2, %r6, bgt_else.9249
"00111111011111100000000000000000",	-- 8947: 	sw	%r27, [%sp + 0]
"00111100011111100000000000000001",	-- 8948: 	sw	%r3, [%sp + 1]
"00111100100111100000000000000010",	-- 8949: 	sw	%r4, [%sp + 2]
"00111100101111100000000000000011",	-- 8950: 	sw	%r5, [%sp + 3]
"00111100010111100000000000000100",	-- 8951: 	sw	%r2, [%sp + 4]
"00111100001111100000000000000101",	-- 8952: 	sw	%r1, [%sp + 5]
"00111111111111100000000000000110",	-- 8953: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8954: 	addi	%sp, %sp, 7
"01011000000000000010000111001011",	-- 8955: 	jal	get_surface_id.2941
"10101011110111100000000000000111",	-- 8956: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8957: 	lw	%ra, [%sp + 6]
"11001100000000100000000000000000",	-- 8958: 	lli	%r2, 0
"00110000010000010000000001010100",	-- 8959: 	bgt	%r2, %r1, bgt_else.9250
"00111011110000010000000000000101",	-- 8960: 	lw	%r1, [%sp + 5]
"00111111111111100000000000000110",	-- 8961: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8962: 	addi	%sp, %sp, 7
"01011000000000000000011010101010",	-- 8963: 	jal	p_calc_diffuse.2670
"10101011110111100000000000000111",	-- 8964: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8965: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000100",	-- 8966: 	lw	%r2, [%sp + 4]
"10000100001000100000100000000000",	-- 8967: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 8968: 	lw	%r1, [%r1 + 0]
"11001100000000110000000000000000",	-- 8969: 	lli	%r3, 0
"00101000001000110000000000000010",	-- 8970: 	bneq	%r1, %r3, bneq_else.9251
"01010100000000000010001101001100",	-- 8971: 	j	bneq_cont.9252
	-- bneq_else.9251:
"00111011110000010000000000000101",	-- 8972: 	lw	%r1, [%sp + 5]
"00111111111111100000000000000110",	-- 8973: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 8974: 	addi	%sp, %sp, 7
"01011000000000000000011010110000",	-- 8975: 	jal	p_group_id.2676
"10101011110111100000000000000111",	-- 8976: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 8977: 	lw	%ra, [%sp + 6]
"00111011110000100000000000000011",	-- 8978: 	lw	%r2, [%sp + 3]
"00111100001111100000000000000110",	-- 8979: 	sw	%r1, [%sp + 6]
"10000100000000100000100000000000",	-- 8980: 	add	%r1, %r0, %r2
"00111111111111100000000000000111",	-- 8981: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 8982: 	addi	%sp, %sp, 8
"01011000000000000000010100111010",	-- 8983: 	jal	vecbzero.2584
"10101011110111100000000000001000",	-- 8984: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8985: 	lw	%ra, [%sp + 7]
"00111011110000010000000000000101",	-- 8986: 	lw	%r1, [%sp + 5]
"00111111111111100000000000000111",	-- 8987: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 8988: 	addi	%sp, %sp, 8
"01011000000000000000011010111010",	-- 8989: 	jal	p_nvectors.2681
"10101011110111100000000000001000",	-- 8990: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 8991: 	lw	%ra, [%sp + 7]
"00111011110000100000000000000101",	-- 8992: 	lw	%r2, [%sp + 5]
"00111100001111100000000000000111",	-- 8993: 	sw	%r1, [%sp + 7]
"10000100000000100000100000000000",	-- 8994: 	add	%r1, %r0, %r2
"00111111111111100000000000001000",	-- 8995: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 8996: 	addi	%sp, %sp, 9
"01011000000000000000011010100110",	-- 8997: 	jal	p_intersection_points.2666
"10101011110111100000000000001001",	-- 8998: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 8999: 	lw	%ra, [%sp + 8]
"00111011110000100000000000000110",	-- 9000: 	lw	%r2, [%sp + 6]
"00111011110000110000000000000010",	-- 9001: 	lw	%r3, [%sp + 2]
"10000100011000100001000000000000",	-- 9002: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 9003: 	lw	%r2, [%r2 + 0]
"00111011110000110000000000000100",	-- 9004: 	lw	%r3, [%sp + 4]
"00111011110001000000000000000111",	-- 9005: 	lw	%r4, [%sp + 7]
"10000100100000110010000000000000",	-- 9006: 	add	%r4, %r4, %r3
"00111000100001000000000000000000",	-- 9007: 	lw	%r4, [%r4 + 0]
"10000100001000110000100000000000",	-- 9008: 	add	%r1, %r1, %r3
"00111000001000010000000000000000",	-- 9009: 	lw	%r1, [%r1 + 0]
"00111011110110110000000000000001",	-- 9010: 	lw	%r27, [%sp + 1]
"10000100000000010001100000000000",	-- 9011: 	add	%r3, %r0, %r1
"10000100000000100000100000000000",	-- 9012: 	add	%r1, %r0, %r2
"10000100000001000001000000000000",	-- 9013: 	add	%r2, %r0, %r4
"00111111111111100000000000001000",	-- 9014: 	sw	%ra, [%sp + 8]
"00111011011110100000000000000000",	-- 9015: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001001",	-- 9016: 	addi	%sp, %sp, 9
"01010011010000000000000000000000",	-- 9017: 	jalr	%r26
"10101011110111100000000000001001",	-- 9018: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 9019: 	lw	%ra, [%sp + 8]
"00111011110000010000000000000101",	-- 9020: 	lw	%r1, [%sp + 5]
"00111111111111100000000000001000",	-- 9021: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 9022: 	addi	%sp, %sp, 9
"01011000000000000000011010101110",	-- 9023: 	jal	p_received_ray_20percent.2674
"10101011110111100000000000001001",	-- 9024: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 9025: 	lw	%ra, [%sp + 8]
"00111011110000100000000000000100",	-- 9026: 	lw	%r2, [%sp + 4]
"10000100001000100000100000000000",	-- 9027: 	add	%r1, %r1, %r2
"00111000001000010000000000000000",	-- 9028: 	lw	%r1, [%r1 + 0]
"00111011110000110000000000000011",	-- 9029: 	lw	%r3, [%sp + 3]
"10000100000000110001000000000000",	-- 9030: 	add	%r2, %r0, %r3
"00111111111111100000000000001000",	-- 9031: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 9032: 	addi	%sp, %sp, 9
"01011000000000000000010100111101",	-- 9033: 	jal	veccpy.2586
"10101011110111100000000000001001",	-- 9034: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 9035: 	lw	%ra, [%sp + 8]
	-- bneq_cont.9252:
"11001100000000010000000000000001",	-- 9036: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 9037: 	lw	%r2, [%sp + 4]
"10000100010000010001000000000000",	-- 9038: 	add	%r2, %r2, %r1
"00111011110000010000000000000101",	-- 9039: 	lw	%r1, [%sp + 5]
"00111011110110110000000000000000",	-- 9040: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 9041: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 9042: 	jr	%r26
	-- bgt_else.9250:
"01001111111000000000000000000000",	-- 9043: 	jr	%ra
	-- bgt_else.9249:
"01001111111000000000000000000000",	-- 9044: 	jr	%ra
	-- pretrace_pixels.2966:
"00111011011001000000000000001001",	-- 9045: 	lw	%r4, [%r27 + 9]
"00111011011001010000000000001000",	-- 9046: 	lw	%r5, [%r27 + 8]
"00111011011001100000000000000111",	-- 9047: 	lw	%r6, [%r27 + 7]
"00111011011001110000000000000110",	-- 9048: 	lw	%r7, [%r27 + 6]
"00111011011010000000000000000101",	-- 9049: 	lw	%r8, [%r27 + 5]
"00111011011010010000000000000100",	-- 9050: 	lw	%r9, [%r27 + 4]
"00111011011010100000000000000011",	-- 9051: 	lw	%r10, [%r27 + 3]
"00111011011010110000000000000010",	-- 9052: 	lw	%r11, [%r27 + 2]
"00111011011011000000000000000001",	-- 9053: 	lw	%r12, [%r27 + 1]
"11001100000011010000000000000000",	-- 9054: 	lli	%r13, 0
"00110001101000100000000010100100",	-- 9055: 	bgt	%r13, %r2, bgt_else.9255
"11001100000011010000000000000000",	-- 9056: 	lli	%r13, 0
"10000101000011010100000000000000",	-- 9057: 	add	%r8, %r8, %r13
"10010001000000110000000000000000",	-- 9058: 	lf	%f3, [%r8 + 0]
"11001100000010000000000000000000",	-- 9059: 	lli	%r8, 0
"10000101100010000100000000000000",	-- 9060: 	add	%r8, %r12, %r8
"00111001000010000000000000000000",	-- 9061: 	lw	%r8, [%r8 + 0]
"10001000010010000100000000000000",	-- 9062: 	sub	%r8, %r2, %r8
"00111111011111100000000000000000",	-- 9063: 	sw	%r27, [%sp + 0]
"00111101011111100000000000000001",	-- 9064: 	sw	%r11, [%sp + 1]
"00111100011111100000000000000010",	-- 9065: 	sw	%r3, [%sp + 2]
"00111100101111100000000000000011",	-- 9066: 	sw	%r5, [%sp + 3]
"00111100010111100000000000000100",	-- 9067: 	sw	%r2, [%sp + 4]
"00111100001111100000000000000101",	-- 9068: 	sw	%r1, [%sp + 5]
"00111100100111100000000000000110",	-- 9069: 	sw	%r4, [%sp + 6]
"00111100110111100000000000000111",	-- 9070: 	sw	%r6, [%sp + 7]
"00111101001111100000000000001000",	-- 9071: 	sw	%r9, [%sp + 8]
"10110000010111100000000000001001",	-- 9072: 	sf	%f2, [%sp + 9]
"10110000001111100000000000001010",	-- 9073: 	sf	%f1, [%sp + 10]
"00111101010111100000000000001011",	-- 9074: 	sw	%r10, [%sp + 11]
"10110000000111100000000000001100",	-- 9075: 	sf	%f0, [%sp + 12]
"00111100111111100000000000001101",	-- 9076: 	sw	%r7, [%sp + 13]
"10110000011111100000000000001110",	-- 9077: 	sf	%f3, [%sp + 14]
"10000100000010000000100000000000",	-- 9078: 	add	%r1, %r0, %r8
"00111111111111100000000000001111",	-- 9079: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9080: 	addi	%sp, %sp, 16
"01011000000000000010101000101100",	-- 9081: 	jal	yj_float_of_int
"10101011110111100000000000010000",	-- 9082: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9083: 	lw	%ra, [%sp + 15]
"10010011110000010000000000001110",	-- 9084: 	lf	%f1, [%sp + 14]
"11101000001000000000000000000000",	-- 9085: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 9086: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 9087: 	lli	%r2, 0
"00111011110000110000000000001101",	-- 9088: 	lw	%r3, [%sp + 13]
"10000100011000100001000000000000",	-- 9089: 	add	%r2, %r3, %r2
"10010000010000010000000000000000",	-- 9090: 	lf	%f1, [%r2 + 0]
"11101000000000010000100000000000",	-- 9091: 	mulf	%f1, %f0, %f1
"10010011110000100000000000001100",	-- 9092: 	lf	%f2, [%sp + 12]
"11100000001000100000100000000000",	-- 9093: 	addf	%f1, %f1, %f2
"00111011110000100000000000001011",	-- 9094: 	lw	%r2, [%sp + 11]
"10000100010000010000100000000000",	-- 9095: 	add	%r1, %r2, %r1
"10110000001000010000000000000000",	-- 9096: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000001",	-- 9097: 	lli	%r1, 1
"11001100000001000000000000000001",	-- 9098: 	lli	%r4, 1
"10000100011001000010000000000000",	-- 9099: 	add	%r4, %r3, %r4
"10010000100000010000000000000000",	-- 9100: 	lf	%f1, [%r4 + 0]
"11101000000000010000100000000000",	-- 9101: 	mulf	%f1, %f0, %f1
"10010011110000110000000000001010",	-- 9102: 	lf	%f3, [%sp + 10]
"11100000001000110000100000000000",	-- 9103: 	addf	%f1, %f1, %f3
"10000100010000010000100000000000",	-- 9104: 	add	%r1, %r2, %r1
"10110000001000010000000000000000",	-- 9105: 	sf	%f1, [%r1 + 0]
"11001100000000010000000000000010",	-- 9106: 	lli	%r1, 2
"11001100000001000000000000000010",	-- 9107: 	lli	%r4, 2
"10000100011001000001100000000000",	-- 9108: 	add	%r3, %r3, %r4
"10010000011000010000000000000000",	-- 9109: 	lf	%f1, [%r3 + 0]
"11101000000000010000000000000000",	-- 9110: 	mulf	%f0, %f0, %f1
"10010011110000010000000000001001",	-- 9111: 	lf	%f1, [%sp + 9]
"11100000000000010000000000000000",	-- 9112: 	addf	%f0, %f0, %f1
"10000100010000010000100000000000",	-- 9113: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 9114: 	sf	%f0, [%r1 + 0]
"11001100000000010000000000000000",	-- 9115: 	lli	%r1, 0
"10000100000000101101000000000000",	-- 9116: 	add	%r26, %r0, %r2
"10000100000000010001000000000000",	-- 9117: 	add	%r2, %r0, %r1
"10000100000110100000100000000000",	-- 9118: 	add	%r1, %r0, %r26
"00111111111111100000000000001111",	-- 9119: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9120: 	addi	%sp, %sp, 16
"01011000000000000000010101010000",	-- 9121: 	jal	vecunit_sgn.2594
"10101011110111100000000000010000",	-- 9122: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9123: 	lw	%ra, [%sp + 15]
"00111011110000010000000000001000",	-- 9124: 	lw	%r1, [%sp + 8]
"00111111111111100000000000001111",	-- 9125: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9126: 	addi	%sp, %sp, 16
"01011000000000000000010100111010",	-- 9127: 	jal	vecbzero.2584
"10101011110111100000000000010000",	-- 9128: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9129: 	lw	%ra, [%sp + 15]
"00111011110000010000000000000111",	-- 9130: 	lw	%r1, [%sp + 7]
"00111011110000100000000000000110",	-- 9131: 	lw	%r2, [%sp + 6]
"00111111111111100000000000001111",	-- 9132: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9133: 	addi	%sp, %sp, 16
"01011000000000000000010100111101",	-- 9134: 	jal	veccpy.2586
"10101011110111100000000000010000",	-- 9135: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9136: 	lw	%ra, [%sp + 15]
"11001100000000010000000000000000",	-- 9137: 	lli	%r1, 0
"00010100000000000000000000000000",	-- 9138: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 9139: 	lhif	%f0, 1.000000
"00111011110000100000000000000100",	-- 9140: 	lw	%r2, [%sp + 4]
"00111011110000110000000000000101",	-- 9141: 	lw	%r3, [%sp + 5]
"10000100011000100010000000000000",	-- 9142: 	add	%r4, %r3, %r2
"00111000100001000000000000000000",	-- 9143: 	lw	%r4, [%r4 + 0]
"00010100000000010000000000000000",	-- 9144: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 9145: 	lhif	%f1, 0.000000
"00111011110001010000000000001011",	-- 9146: 	lw	%r5, [%sp + 11]
"00111011110110110000000000000011",	-- 9147: 	lw	%r27, [%sp + 3]
"10000100000001000001100000000000",	-- 9148: 	add	%r3, %r0, %r4
"10000100000001010001000000000000",	-- 9149: 	add	%r2, %r0, %r5
"00111111111111100000000000001111",	-- 9150: 	sw	%ra, [%sp + 15]
"00111011011110100000000000000000",	-- 9151: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010000",	-- 9152: 	addi	%sp, %sp, 16
"01010011010000000000000000000000",	-- 9153: 	jalr	%r26
"10101011110111100000000000010000",	-- 9154: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9155: 	lw	%ra, [%sp + 15]
"00111011110000010000000000000100",	-- 9156: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000101",	-- 9157: 	lw	%r2, [%sp + 5]
"10000100010000010001100000000000",	-- 9158: 	add	%r3, %r2, %r1
"00111000011000110000000000000000",	-- 9159: 	lw	%r3, [%r3 + 0]
"10000100000000110000100000000000",	-- 9160: 	add	%r1, %r0, %r3
"00111111111111100000000000001111",	-- 9161: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9162: 	addi	%sp, %sp, 16
"01011000000000000000011010100100",	-- 9163: 	jal	p_rgb.2664
"10101011110111100000000000010000",	-- 9164: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9165: 	lw	%ra, [%sp + 15]
"00111011110000100000000000001000",	-- 9166: 	lw	%r2, [%sp + 8]
"00111111111111100000000000001111",	-- 9167: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9168: 	addi	%sp, %sp, 16
"01011000000000000000010100111101",	-- 9169: 	jal	veccpy.2586
"10101011110111100000000000010000",	-- 9170: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9171: 	lw	%ra, [%sp + 15]
"00111011110000010000000000000100",	-- 9172: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000101",	-- 9173: 	lw	%r2, [%sp + 5]
"10000100010000010001100000000000",	-- 9174: 	add	%r3, %r2, %r1
"00111000011000110000000000000000",	-- 9175: 	lw	%r3, [%r3 + 0]
"00111011110001000000000000000010",	-- 9176: 	lw	%r4, [%sp + 2]
"10000100000001000001000000000000",	-- 9177: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 9178: 	add	%r1, %r0, %r3
"00111111111111100000000000001111",	-- 9179: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9180: 	addi	%sp, %sp, 16
"01011000000000000000011010110101",	-- 9181: 	jal	p_set_group_id.2678
"10101011110111100000000000010000",	-- 9182: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9183: 	lw	%ra, [%sp + 15]
"00111011110000010000000000000100",	-- 9184: 	lw	%r1, [%sp + 4]
"00111011110000100000000000000101",	-- 9185: 	lw	%r2, [%sp + 5]
"10000100010000010001100000000000",	-- 9186: 	add	%r3, %r2, %r1
"00111000011000110000000000000000",	-- 9187: 	lw	%r3, [%r3 + 0]
"11001100000001000000000000000000",	-- 9188: 	lli	%r4, 0
"00111011110110110000000000000001",	-- 9189: 	lw	%r27, [%sp + 1]
"10000100000001000001000000000000",	-- 9190: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 9191: 	add	%r1, %r0, %r3
"00111111111111100000000000001111",	-- 9192: 	sw	%ra, [%sp + 15]
"00111011011110100000000000000000",	-- 9193: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010000",	-- 9194: 	addi	%sp, %sp, 16
"01010011010000000000000000000000",	-- 9195: 	jalr	%r26
"10101011110111100000000000010000",	-- 9196: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9197: 	lw	%ra, [%sp + 15]
"11001100000000010000000000000001",	-- 9198: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 9199: 	lw	%r2, [%sp + 4]
"10001000010000010000100000000000",	-- 9200: 	sub	%r1, %r2, %r1
"11001100000000100000000000000001",	-- 9201: 	lli	%r2, 1
"00111011110000110000000000000010",	-- 9202: 	lw	%r3, [%sp + 2]
"00111100001111100000000000001111",	-- 9203: 	sw	%r1, [%sp + 15]
"10000100000000110000100000000000",	-- 9204: 	add	%r1, %r0, %r3
"00111111111111100000000000010000",	-- 9205: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 9206: 	addi	%sp, %sp, 17
"01011000000000000000010100011111",	-- 9207: 	jal	add_mod5.2573
"10101011110111100000000000010001",	-- 9208: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 9209: 	lw	%ra, [%sp + 16]
"10000100000000010001100000000000",	-- 9210: 	add	%r3, %r0, %r1
"10010011110000000000000000001100",	-- 9211: 	lf	%f0, [%sp + 12]
"10010011110000010000000000001010",	-- 9212: 	lf	%f1, [%sp + 10]
"10010011110000100000000000001001",	-- 9213: 	lf	%f2, [%sp + 9]
"00111011110000010000000000000101",	-- 9214: 	lw	%r1, [%sp + 5]
"00111011110000100000000000001111",	-- 9215: 	lw	%r2, [%sp + 15]
"00111011110110110000000000000000",	-- 9216: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 9217: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 9218: 	jr	%r26
	-- bgt_else.9255:
"01001111111000000000000000000000",	-- 9219: 	jr	%ra
	-- pretrace_line.2973:
"00111011011001000000000000000110",	-- 9220: 	lw	%r4, [%r27 + 6]
"00111011011001010000000000000101",	-- 9221: 	lw	%r5, [%r27 + 5]
"00111011011001100000000000000100",	-- 9222: 	lw	%r6, [%r27 + 4]
"00111011011001110000000000000011",	-- 9223: 	lw	%r7, [%r27 + 3]
"00111011011010000000000000000010",	-- 9224: 	lw	%r8, [%r27 + 2]
"00111011011010010000000000000001",	-- 9225: 	lw	%r9, [%r27 + 1]
"11001100000010100000000000000000",	-- 9226: 	lli	%r10, 0
"10000100110010100011000000000000",	-- 9227: 	add	%r6, %r6, %r10
"10010000110000000000000000000000",	-- 9228: 	lf	%f0, [%r6 + 0]
"11001100000001100000000000000001",	-- 9229: 	lli	%r6, 1
"10000101001001100011000000000000",	-- 9230: 	add	%r6, %r9, %r6
"00111000110001100000000000000000",	-- 9231: 	lw	%r6, [%r6 + 0]
"10001000010001100001000000000000",	-- 9232: 	sub	%r2, %r2, %r6
"00111100011111100000000000000000",	-- 9233: 	sw	%r3, [%sp + 0]
"00111100001111100000000000000001",	-- 9234: 	sw	%r1, [%sp + 1]
"00111100111111100000000000000010",	-- 9235: 	sw	%r7, [%sp + 2]
"00111101000111100000000000000011",	-- 9236: 	sw	%r8, [%sp + 3]
"00111100100111100000000000000100",	-- 9237: 	sw	%r4, [%sp + 4]
"00111100101111100000000000000101",	-- 9238: 	sw	%r5, [%sp + 5]
"10110000000111100000000000000110",	-- 9239: 	sf	%f0, [%sp + 6]
"10000100000000100000100000000000",	-- 9240: 	add	%r1, %r0, %r2
"00111111111111100000000000000111",	-- 9241: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 9242: 	addi	%sp, %sp, 8
"01011000000000000010101000101100",	-- 9243: 	jal	yj_float_of_int
"10101011110111100000000000001000",	-- 9244: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 9245: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000110",	-- 9246: 	lf	%f1, [%sp + 6]
"11101000001000000000000000000000",	-- 9247: 	mulf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 9248: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 9249: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 9250: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 9251: 	lf	%f1, [%r1 + 0]
"11101000000000010000100000000000",	-- 9252: 	mulf	%f1, %f0, %f1
"11001100000000010000000000000000",	-- 9253: 	lli	%r1, 0
"00111011110000110000000000000100",	-- 9254: 	lw	%r3, [%sp + 4]
"10000100011000010000100000000000",	-- 9255: 	add	%r1, %r3, %r1
"10010000001000100000000000000000",	-- 9256: 	lf	%f2, [%r1 + 0]
"11100000001000100000100000000000",	-- 9257: 	addf	%f1, %f1, %f2
"11001100000000010000000000000001",	-- 9258: 	lli	%r1, 1
"10000100010000010000100000000000",	-- 9259: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 9260: 	lf	%f2, [%r1 + 0]
"11101000000000100001000000000000",	-- 9261: 	mulf	%f2, %f0, %f2
"11001100000000010000000000000001",	-- 9262: 	lli	%r1, 1
"10000100011000010000100000000000",	-- 9263: 	add	%r1, %r3, %r1
"10010000001000110000000000000000",	-- 9264: 	lf	%f3, [%r1 + 0]
"11100000010000110001000000000000",	-- 9265: 	addf	%f2, %f2, %f3
"11001100000000010000000000000010",	-- 9266: 	lli	%r1, 2
"10000100010000010000100000000000",	-- 9267: 	add	%r1, %r2, %r1
"10010000001000110000000000000000",	-- 9268: 	lf	%f3, [%r1 + 0]
"11101000000000110000000000000000",	-- 9269: 	mulf	%f0, %f0, %f3
"11001100000000010000000000000010",	-- 9270: 	lli	%r1, 2
"10000100011000010000100000000000",	-- 9271: 	add	%r1, %r3, %r1
"10010000001000110000000000000000",	-- 9272: 	lf	%f3, [%r1 + 0]
"11100000000000110000000000000000",	-- 9273: 	addf	%f0, %f0, %f3
"11001100000000010000000000000000",	-- 9274: 	lli	%r1, 0
"00111011110000100000000000000011",	-- 9275: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 9276: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 9277: 	lw	%r1, [%r1 + 0]
"11001100000000100000000000000001",	-- 9278: 	lli	%r2, 1
"10001000001000100001000000000000",	-- 9279: 	sub	%r2, %r1, %r2
"00111011110000010000000000000001",	-- 9280: 	lw	%r1, [%sp + 1]
"00111011110000110000000000000000",	-- 9281: 	lw	%r3, [%sp + 0]
"00111011110110110000000000000010",	-- 9282: 	lw	%r27, [%sp + 2]
"00001100010111110000000000000000",	-- 9283: 	movf	%f31, %f2
"00001100000000100000000000000000",	-- 9284: 	movf	%f2, %f0
"00001100001000000000000000000000",	-- 9285: 	movf	%f0, %f1
"00001111111000010000000000000000",	-- 9286: 	movf	%f1, %f31
"00111011011110100000000000000000",	-- 9287: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 9288: 	jr	%r26
	-- scan_pixel.2977:
"00111011011001100000000000000110",	-- 9289: 	lw	%r6, [%r27 + 6]
"00111011011001110000000000000101",	-- 9290: 	lw	%r7, [%r27 + 5]
"00111011011010000000000000000100",	-- 9291: 	lw	%r8, [%r27 + 4]
"00111011011010010000000000000011",	-- 9292: 	lw	%r9, [%r27 + 3]
"00111011011010100000000000000010",	-- 9293: 	lw	%r10, [%r27 + 2]
"00111011011010110000000000000001",	-- 9294: 	lw	%r11, [%r27 + 1]
"11001100000011000000000000000000",	-- 9295: 	lli	%r12, 0
"10000101010011000101000000000000",	-- 9296: 	add	%r10, %r10, %r12
"00111001010010100000000000000000",	-- 9297: 	lw	%r10, [%r10 + 0]
"00110001010000010000000000000010",	-- 9298: 	bgt	%r10, %r1, bgt_else.9257
"01001111111000000000000000000000",	-- 9299: 	jr	%ra
	-- bgt_else.9257:
"10000100100000010101000000000000",	-- 9300: 	add	%r10, %r4, %r1
"00111001010010100000000000000000",	-- 9301: 	lw	%r10, [%r10 + 0]
"00111111011111100000000000000000",	-- 9302: 	sw	%r27, [%sp + 0]
"00111100110111100000000000000001",	-- 9303: 	sw	%r6, [%sp + 1]
"00111100011111100000000000000010",	-- 9304: 	sw	%r3, [%sp + 2]
"00111100111111100000000000000011",	-- 9305: 	sw	%r7, [%sp + 3]
"00111101011111100000000000000100",	-- 9306: 	sw	%r11, [%sp + 4]
"00111100100111100000000000000101",	-- 9307: 	sw	%r4, [%sp + 5]
"00111100101111100000000000000110",	-- 9308: 	sw	%r5, [%sp + 6]
"00111100010111100000000000000111",	-- 9309: 	sw	%r2, [%sp + 7]
"00111100001111100000000000001000",	-- 9310: 	sw	%r1, [%sp + 8]
"00111101001111100000000000001001",	-- 9311: 	sw	%r9, [%sp + 9]
"00111101000111100000000000001010",	-- 9312: 	sw	%r8, [%sp + 10]
"10000100000010100000100000000000",	-- 9313: 	add	%r1, %r0, %r10
"00111111111111100000000000001011",	-- 9314: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 9315: 	addi	%sp, %sp, 12
"01011000000000000000011010100100",	-- 9316: 	jal	p_rgb.2664
"10101011110111100000000000001100",	-- 9317: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9318: 	lw	%ra, [%sp + 11]
"10000100000000010001000000000000",	-- 9319: 	add	%r2, %r0, %r1
"00111011110000010000000000001010",	-- 9320: 	lw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 9321: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 9322: 	addi	%sp, %sp, 12
"01011000000000000000010100111101",	-- 9323: 	jal	veccpy.2586
"10101011110111100000000000001100",	-- 9324: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9325: 	lw	%ra, [%sp + 11]
"00111011110000010000000000001000",	-- 9326: 	lw	%r1, [%sp + 8]
"00111011110000100000000000000111",	-- 9327: 	lw	%r2, [%sp + 7]
"00111011110000110000000000000110",	-- 9328: 	lw	%r3, [%sp + 6]
"00111011110110110000000000001001",	-- 9329: 	lw	%r27, [%sp + 9]
"00111111111111100000000000001011",	-- 9330: 	sw	%ra, [%sp + 11]
"00111011011110100000000000000000",	-- 9331: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001100",	-- 9332: 	addi	%sp, %sp, 12
"01010011010000000000000000000000",	-- 9333: 	jalr	%r26
"10101011110111100000000000001100",	-- 9334: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9335: 	lw	%ra, [%sp + 11]
"11001100000000100000000000000000",	-- 9336: 	lli	%r2, 0
"00101000001000100000000000010000",	-- 9337: 	bneq	%r1, %r2, bneq_else.9259
"00111011110000010000000000001000",	-- 9338: 	lw	%r1, [%sp + 8]
"00111011110000100000000000000101",	-- 9339: 	lw	%r2, [%sp + 5]
"10000100010000010001100000000000",	-- 9340: 	add	%r3, %r2, %r1
"00111000011000110000000000000000",	-- 9341: 	lw	%r3, [%r3 + 0]
"11001100000001000000000000000000",	-- 9342: 	lli	%r4, 0
"00111011110110110000000000000100",	-- 9343: 	lw	%r27, [%sp + 4]
"10000100000001000001000000000000",	-- 9344: 	add	%r2, %r0, %r4
"10000100000000110000100000000000",	-- 9345: 	add	%r1, %r0, %r3
"00111111111111100000000000001011",	-- 9346: 	sw	%ra, [%sp + 11]
"00111011011110100000000000000000",	-- 9347: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001100",	-- 9348: 	addi	%sp, %sp, 12
"01010011010000000000000000000000",	-- 9349: 	jalr	%r26
"10101011110111100000000000001100",	-- 9350: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9351: 	lw	%ra, [%sp + 11]
"01010100000000000010010010010110",	-- 9352: 	j	bneq_cont.9260
	-- bneq_else.9259:
"11001100000001100000000000000000",	-- 9353: 	lli	%r6, 0
"00111011110000010000000000001000",	-- 9354: 	lw	%r1, [%sp + 8]
"00111011110000100000000000000111",	-- 9355: 	lw	%r2, [%sp + 7]
"00111011110000110000000000000010",	-- 9356: 	lw	%r3, [%sp + 2]
"00111011110001000000000000000101",	-- 9357: 	lw	%r4, [%sp + 5]
"00111011110001010000000000000110",	-- 9358: 	lw	%r5, [%sp + 6]
"00111011110110110000000000000011",	-- 9359: 	lw	%r27, [%sp + 3]
"00111111111111100000000000001011",	-- 9360: 	sw	%ra, [%sp + 11]
"00111011011110100000000000000000",	-- 9361: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001100",	-- 9362: 	addi	%sp, %sp, 12
"01010011010000000000000000000000",	-- 9363: 	jalr	%r26
"10101011110111100000000000001100",	-- 9364: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9365: 	lw	%ra, [%sp + 11]
	-- bneq_cont.9260:
"00111011110110110000000000000001",	-- 9366: 	lw	%r27, [%sp + 1]
"00111111111111100000000000001011",	-- 9367: 	sw	%ra, [%sp + 11]
"00111011011110100000000000000000",	-- 9368: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001100",	-- 9369: 	addi	%sp, %sp, 12
"01010011010000000000000000000000",	-- 9370: 	jalr	%r26
"10101011110111100000000000001100",	-- 9371: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9372: 	lw	%ra, [%sp + 11]
"11001100000000010000000000000001",	-- 9373: 	lli	%r1, 1
"00111011110000100000000000001000",	-- 9374: 	lw	%r2, [%sp + 8]
"10000100010000010000100000000000",	-- 9375: 	add	%r1, %r2, %r1
"00111011110000100000000000000111",	-- 9376: 	lw	%r2, [%sp + 7]
"00111011110000110000000000000010",	-- 9377: 	lw	%r3, [%sp + 2]
"00111011110001000000000000000101",	-- 9378: 	lw	%r4, [%sp + 5]
"00111011110001010000000000000110",	-- 9379: 	lw	%r5, [%sp + 6]
"00111011110110110000000000000000",	-- 9380: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 9381: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 9382: 	jr	%r26
	-- scan_line.2983:
"00111011011001100000000000000011",	-- 9383: 	lw	%r6, [%r27 + 3]
"00111011011001110000000000000010",	-- 9384: 	lw	%r7, [%r27 + 2]
"00111011011010000000000000000001",	-- 9385: 	lw	%r8, [%r27 + 1]
"11001100000010010000000000000001",	-- 9386: 	lli	%r9, 1
"10000101000010010100100000000000",	-- 9387: 	add	%r9, %r8, %r9
"00111001001010010000000000000000",	-- 9388: 	lw	%r9, [%r9 + 0]
"00110001001000010000000000000010",	-- 9389: 	bgt	%r9, %r1, bgt_else.9261
"01001111111000000000000000000000",	-- 9390: 	jr	%ra
	-- bgt_else.9261:
"11001100000010010000000000000001",	-- 9391: 	lli	%r9, 1
"10000101000010010100000000000000",	-- 9392: 	add	%r8, %r8, %r9
"00111001000010000000000000000000",	-- 9393: 	lw	%r8, [%r8 + 0]
"11001100000010010000000000000001",	-- 9394: 	lli	%r9, 1
"10001001000010010100000000000000",	-- 9395: 	sub	%r8, %r8, %r9
"00111111011111100000000000000000",	-- 9396: 	sw	%r27, [%sp + 0]
"00111100101111100000000000000001",	-- 9397: 	sw	%r5, [%sp + 1]
"00111100100111100000000000000010",	-- 9398: 	sw	%r4, [%sp + 2]
"00111100011111100000000000000011",	-- 9399: 	sw	%r3, [%sp + 3]
"00111100010111100000000000000100",	-- 9400: 	sw	%r2, [%sp + 4]
"00111100001111100000000000000101",	-- 9401: 	sw	%r1, [%sp + 5]
"00111100110111100000000000000110",	-- 9402: 	sw	%r6, [%sp + 6]
"00110001000000010000000000000010",	-- 9403: 	bgt	%r8, %r1, bgt_else.9263
"01010100000000000010010011001001",	-- 9404: 	j	bgt_cont.9264
	-- bgt_else.9263:
"11001100000010000000000000000001",	-- 9405: 	lli	%r8, 1
"10000100001010000100000000000000",	-- 9406: 	add	%r8, %r1, %r8
"10000100000001010001100000000000",	-- 9407: 	add	%r3, %r0, %r5
"10000100000010000001000000000000",	-- 9408: 	add	%r2, %r0, %r8
"10000100000001000000100000000000",	-- 9409: 	add	%r1, %r0, %r4
"10000100000001111101100000000000",	-- 9410: 	add	%r27, %r0, %r7
"00111111111111100000000000000111",	-- 9411: 	sw	%ra, [%sp + 7]
"00111011011110100000000000000000",	-- 9412: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001000",	-- 9413: 	addi	%sp, %sp, 8
"01010011010000000000000000000000",	-- 9414: 	jalr	%r26
"10101011110111100000000000001000",	-- 9415: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 9416: 	lw	%ra, [%sp + 7]
	-- bgt_cont.9264:
"11001100000000010000000000000000",	-- 9417: 	lli	%r1, 0
"00111011110000100000000000000101",	-- 9418: 	lw	%r2, [%sp + 5]
"00111011110000110000000000000100",	-- 9419: 	lw	%r3, [%sp + 4]
"00111011110001000000000000000011",	-- 9420: 	lw	%r4, [%sp + 3]
"00111011110001010000000000000010",	-- 9421: 	lw	%r5, [%sp + 2]
"00111011110110110000000000000110",	-- 9422: 	lw	%r27, [%sp + 6]
"00111111111111100000000000000111",	-- 9423: 	sw	%ra, [%sp + 7]
"00111011011110100000000000000000",	-- 9424: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001000",	-- 9425: 	addi	%sp, %sp, 8
"01010011010000000000000000000000",	-- 9426: 	jalr	%r26
"10101011110111100000000000001000",	-- 9427: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 9428: 	lw	%ra, [%sp + 7]
"11001100000000010000000000000001",	-- 9429: 	lli	%r1, 1
"00111011110000100000000000000101",	-- 9430: 	lw	%r2, [%sp + 5]
"10000100010000010000100000000000",	-- 9431: 	add	%r1, %r2, %r1
"11001100000000100000000000000010",	-- 9432: 	lli	%r2, 2
"00111011110000110000000000000001",	-- 9433: 	lw	%r3, [%sp + 1]
"00111100001111100000000000000111",	-- 9434: 	sw	%r1, [%sp + 7]
"10000100000000110000100000000000",	-- 9435: 	add	%r1, %r0, %r3
"00111111111111100000000000001000",	-- 9436: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 9437: 	addi	%sp, %sp, 9
"01011000000000000000010100011111",	-- 9438: 	jal	add_mod5.2573
"10101011110111100000000000001001",	-- 9439: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 9440: 	lw	%ra, [%sp + 8]
"10000100000000010010100000000000",	-- 9441: 	add	%r5, %r0, %r1
"00111011110000010000000000000111",	-- 9442: 	lw	%r1, [%sp + 7]
"00111011110000100000000000000011",	-- 9443: 	lw	%r2, [%sp + 3]
"00111011110000110000000000000010",	-- 9444: 	lw	%r3, [%sp + 2]
"00111011110001000000000000000100",	-- 9445: 	lw	%r4, [%sp + 4]
"00111011110110110000000000000000",	-- 9446: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 9447: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 9448: 	jr	%r26
	-- create_float5x3array.2989:
"11001100000000010000000000000011",	-- 9449: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 9450: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9451: 	lhif	%f0, 0.000000
"00111111111111100000000000000000",	-- 9452: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 9453: 	addi	%sp, %sp, 1
"01011000000000000010101000100100",	-- 9454: 	jal	yj_create_float_array
"10101011110111100000000000000001",	-- 9455: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 9456: 	lw	%ra, [%sp + 0]
"10000100000000010001000000000000",	-- 9457: 	add	%r2, %r0, %r1
"11001100000000010000000000000101",	-- 9458: 	lli	%r1, 5
"00111111111111100000000000000000",	-- 9459: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 9460: 	addi	%sp, %sp, 1
"01011000000000000010101000011100",	-- 9461: 	jal	yj_create_array
"10101011110111100000000000000001",	-- 9462: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 9463: 	lw	%ra, [%sp + 0]
"11001100000000100000000000000001",	-- 9464: 	lli	%r2, 1
"11001100000000110000000000000011",	-- 9465: 	lli	%r3, 3
"00010100000000000000000000000000",	-- 9466: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9467: 	lhif	%f0, 0.000000
"00111100010111100000000000000000",	-- 9468: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 9469: 	sw	%r1, [%sp + 1]
"10000100000000110000100000000000",	-- 9470: 	add	%r1, %r0, %r3
"00111111111111100000000000000010",	-- 9471: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9472: 	addi	%sp, %sp, 3
"01011000000000000010101000100100",	-- 9473: 	jal	yj_create_float_array
"10101011110111100000000000000011",	-- 9474: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9475: 	lw	%ra, [%sp + 2]
"00111011110000100000000000000000",	-- 9476: 	lw	%r2, [%sp + 0]
"00111011110000110000000000000001",	-- 9477: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 9478: 	add	%r2, %r3, %r2
"00111100001000100000000000000000",	-- 9479: 	sw	%r1, [%r2 + 0]
"11001100000000010000000000000010",	-- 9480: 	lli	%r1, 2
"11001100000000100000000000000011",	-- 9481: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 9482: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9483: 	lhif	%f0, 0.000000
"00111100001111100000000000000010",	-- 9484: 	sw	%r1, [%sp + 2]
"10000100000000100000100000000000",	-- 9485: 	add	%r1, %r0, %r2
"00111111111111100000000000000011",	-- 9486: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 9487: 	addi	%sp, %sp, 4
"01011000000000000010101000100100",	-- 9488: 	jal	yj_create_float_array
"10101011110111100000000000000100",	-- 9489: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 9490: 	lw	%ra, [%sp + 3]
"00111011110000100000000000000010",	-- 9491: 	lw	%r2, [%sp + 2]
"00111011110000110000000000000001",	-- 9492: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 9493: 	add	%r2, %r3, %r2
"00111100001000100000000000000000",	-- 9494: 	sw	%r1, [%r2 + 0]
"11001100000000010000000000000011",	-- 9495: 	lli	%r1, 3
"11001100000000100000000000000011",	-- 9496: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 9497: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9498: 	lhif	%f0, 0.000000
"00111100001111100000000000000011",	-- 9499: 	sw	%r1, [%sp + 3]
"10000100000000100000100000000000",	-- 9500: 	add	%r1, %r0, %r2
"00111111111111100000000000000100",	-- 9501: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 9502: 	addi	%sp, %sp, 5
"01011000000000000010101000100100",	-- 9503: 	jal	yj_create_float_array
"10101011110111100000000000000101",	-- 9504: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 9505: 	lw	%ra, [%sp + 4]
"00111011110000100000000000000011",	-- 9506: 	lw	%r2, [%sp + 3]
"00111011110000110000000000000001",	-- 9507: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 9508: 	add	%r2, %r3, %r2
"00111100001000100000000000000000",	-- 9509: 	sw	%r1, [%r2 + 0]
"11001100000000010000000000000100",	-- 9510: 	lli	%r1, 4
"11001100000000100000000000000011",	-- 9511: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 9512: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9513: 	lhif	%f0, 0.000000
"00111100001111100000000000000100",	-- 9514: 	sw	%r1, [%sp + 4]
"10000100000000100000100000000000",	-- 9515: 	add	%r1, %r0, %r2
"00111111111111100000000000000101",	-- 9516: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 9517: 	addi	%sp, %sp, 6
"01011000000000000010101000100100",	-- 9518: 	jal	yj_create_float_array
"10101011110111100000000000000110",	-- 9519: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 9520: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000100",	-- 9521: 	lw	%r2, [%sp + 4]
"00111011110000110000000000000001",	-- 9522: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 9523: 	add	%r2, %r3, %r2
"00111100001000100000000000000000",	-- 9524: 	sw	%r1, [%r2 + 0]
"10000100000000110000100000000000",	-- 9525: 	add	%r1, %r0, %r3
"01001111111000000000000000000000",	-- 9526: 	jr	%ra
	-- create_pixel.2991:
"11001100000000010000000000000011",	-- 9527: 	lli	%r1, 3
"00010100000000000000000000000000",	-- 9528: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9529: 	lhif	%f0, 0.000000
"00111111111111100000000000000000",	-- 9530: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 9531: 	addi	%sp, %sp, 1
"01011000000000000010101000100100",	-- 9532: 	jal	yj_create_float_array
"10101011110111100000000000000001",	-- 9533: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 9534: 	lw	%ra, [%sp + 0]
"00111100001111100000000000000000",	-- 9535: 	sw	%r1, [%sp + 0]
"00111111111111100000000000000001",	-- 9536: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 9537: 	addi	%sp, %sp, 2
"01011000000000000010010011101001",	-- 9538: 	jal	create_float5x3array.2989
"10101011110111100000000000000010",	-- 9539: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 9540: 	lw	%ra, [%sp + 1]
"11001100000000100000000000000101",	-- 9541: 	lli	%r2, 5
"11001100000000110000000000000000",	-- 9542: 	lli	%r3, 0
"00111100001111100000000000000001",	-- 9543: 	sw	%r1, [%sp + 1]
"10000100000000100000100000000000",	-- 9544: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 9545: 	add	%r2, %r0, %r3
"00111111111111100000000000000010",	-- 9546: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9547: 	addi	%sp, %sp, 3
"01011000000000000010101000011100",	-- 9548: 	jal	yj_create_array
"10101011110111100000000000000011",	-- 9549: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9550: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000101",	-- 9551: 	lli	%r2, 5
"11001100000000110000000000000000",	-- 9552: 	lli	%r3, 0
"00111100001111100000000000000010",	-- 9553: 	sw	%r1, [%sp + 2]
"10000100000000100000100000000000",	-- 9554: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 9555: 	add	%r2, %r0, %r3
"00111111111111100000000000000011",	-- 9556: 	sw	%ra, [%sp + 3]
"10100111110111100000000000000100",	-- 9557: 	addi	%sp, %sp, 4
"01011000000000000010101000011100",	-- 9558: 	jal	yj_create_array
"10101011110111100000000000000100",	-- 9559: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 9560: 	lw	%ra, [%sp + 3]
"00111100001111100000000000000011",	-- 9561: 	sw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 9562: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 9563: 	addi	%sp, %sp, 5
"01011000000000000010010011101001",	-- 9564: 	jal	create_float5x3array.2989
"10101011110111100000000000000101",	-- 9565: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 9566: 	lw	%ra, [%sp + 4]
"00111100001111100000000000000100",	-- 9567: 	sw	%r1, [%sp + 4]
"00111111111111100000000000000101",	-- 9568: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 9569: 	addi	%sp, %sp, 6
"01011000000000000010010011101001",	-- 9570: 	jal	create_float5x3array.2989
"10101011110111100000000000000110",	-- 9571: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 9572: 	lw	%ra, [%sp + 5]
"11001100000000100000000000000001",	-- 9573: 	lli	%r2, 1
"11001100000000110000000000000000",	-- 9574: 	lli	%r3, 0
"00111100001111100000000000000101",	-- 9575: 	sw	%r1, [%sp + 5]
"10000100000000100000100000000000",	-- 9576: 	add	%r1, %r0, %r2
"10000100000000110001000000000000",	-- 9577: 	add	%r2, %r0, %r3
"00111111111111100000000000000110",	-- 9578: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 9579: 	addi	%sp, %sp, 7
"01011000000000000010101000011100",	-- 9580: 	jal	yj_create_array
"10101011110111100000000000000111",	-- 9581: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 9582: 	lw	%ra, [%sp + 6]
"00111100001111100000000000000110",	-- 9583: 	sw	%r1, [%sp + 6]
"00111111111111100000000000000111",	-- 9584: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 9585: 	addi	%sp, %sp, 8
"01011000000000000010010011101001",	-- 9586: 	jal	create_float5x3array.2989
"10101011110111100000000000001000",	-- 9587: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 9588: 	lw	%ra, [%sp + 7]
"10000100000111010001000000000000",	-- 9589: 	add	%r2, %r0, %hp
"10100111101111010000000000001000",	-- 9590: 	addi	%hp, %hp, 8
"00111100001000100000000000000111",	-- 9591: 	sw	%r1, [%r2 + 7]
"00111011110000010000000000000110",	-- 9592: 	lw	%r1, [%sp + 6]
"00111100001000100000000000000110",	-- 9593: 	sw	%r1, [%r2 + 6]
"00111011110000010000000000000101",	-- 9594: 	lw	%r1, [%sp + 5]
"00111100001000100000000000000101",	-- 9595: 	sw	%r1, [%r2 + 5]
"00111011110000010000000000000100",	-- 9596: 	lw	%r1, [%sp + 4]
"00111100001000100000000000000100",	-- 9597: 	sw	%r1, [%r2 + 4]
"00111011110000010000000000000011",	-- 9598: 	lw	%r1, [%sp + 3]
"00111100001000100000000000000011",	-- 9599: 	sw	%r1, [%r2 + 3]
"00111011110000010000000000000010",	-- 9600: 	lw	%r1, [%sp + 2]
"00111100001000100000000000000010",	-- 9601: 	sw	%r1, [%r2 + 2]
"00111011110000010000000000000001",	-- 9602: 	lw	%r1, [%sp + 1]
"00111100001000100000000000000001",	-- 9603: 	sw	%r1, [%r2 + 1]
"00111011110000010000000000000000",	-- 9604: 	lw	%r1, [%sp + 0]
"00111100001000100000000000000000",	-- 9605: 	sw	%r1, [%r2 + 0]
"10000100000000100000100000000000",	-- 9606: 	add	%r1, %r0, %r2
"01001111111000000000000000000000",	-- 9607: 	jr	%ra
	-- init_line_elements.2993:
"11001100000000110000000000000000",	-- 9608: 	lli	%r3, 0
"00110000011000100000000000010000",	-- 9609: 	bgt	%r3, %r2, bgt_else.9265
"00111100010111100000000000000000",	-- 9610: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 9611: 	sw	%r1, [%sp + 1]
"00111111111111100000000000000010",	-- 9612: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9613: 	addi	%sp, %sp, 3
"01011000000000000010010100110111",	-- 9614: 	jal	create_pixel.2991
"10101011110111100000000000000011",	-- 9615: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9616: 	lw	%ra, [%sp + 2]
"00111011110000100000000000000000",	-- 9617: 	lw	%r2, [%sp + 0]
"00111011110000110000000000000001",	-- 9618: 	lw	%r3, [%sp + 1]
"10000100011000100010000000000000",	-- 9619: 	add	%r4, %r3, %r2
"00111100001001000000000000000000",	-- 9620: 	sw	%r1, [%r4 + 0]
"11001100000000010000000000000001",	-- 9621: 	lli	%r1, 1
"10001000010000010001000000000000",	-- 9622: 	sub	%r2, %r2, %r1
"10000100000000110000100000000000",	-- 9623: 	add	%r1, %r0, %r3
"01010100000000000010010110001000",	-- 9624: 	j	init_line_elements.2993
	-- bgt_else.9265:
"01001111111000000000000000000000",	-- 9625: 	jr	%ra
	-- create_pixelline.2996:
"00111011011000010000000000000001",	-- 9626: 	lw	%r1, [%r27 + 1]
"11001100000000100000000000000000",	-- 9627: 	lli	%r2, 0
"10000100001000100001000000000000",	-- 9628: 	add	%r2, %r1, %r2
"00111000010000100000000000000000",	-- 9629: 	lw	%r2, [%r2 + 0]
"00111100001111100000000000000000",	-- 9630: 	sw	%r1, [%sp + 0]
"00111100010111100000000000000001",	-- 9631: 	sw	%r2, [%sp + 1]
"00111111111111100000000000000010",	-- 9632: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9633: 	addi	%sp, %sp, 3
"01011000000000000010010100110111",	-- 9634: 	jal	create_pixel.2991
"10101011110111100000000000000011",	-- 9635: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9636: 	lw	%ra, [%sp + 2]
"10000100000000010001000000000000",	-- 9637: 	add	%r2, %r0, %r1
"00111011110000010000000000000001",	-- 9638: 	lw	%r1, [%sp + 1]
"00111111111111100000000000000010",	-- 9639: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9640: 	addi	%sp, %sp, 3
"01011000000000000010101000011100",	-- 9641: 	jal	yj_create_array
"10101011110111100000000000000011",	-- 9642: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9643: 	lw	%ra, [%sp + 2]
"11001100000000100000000000000000",	-- 9644: 	lli	%r2, 0
"00111011110000110000000000000000",	-- 9645: 	lw	%r3, [%sp + 0]
"10000100011000100001000000000000",	-- 9646: 	add	%r2, %r3, %r2
"00111000010000100000000000000000",	-- 9647: 	lw	%r2, [%r2 + 0]
"11001100000000110000000000000010",	-- 9648: 	lli	%r3, 2
"10001000010000110001000000000000",	-- 9649: 	sub	%r2, %r2, %r3
"01010100000000000010010110001000",	-- 9650: 	j	init_line_elements.2993
	-- tan.2998:
"10110000000111100000000000000000",	-- 9651: 	sf	%f0, [%sp + 0]
"00111111111111100000000000000001",	-- 9652: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 9653: 	addi	%sp, %sp, 2
"01011000000000000000010001011001",	-- 9654: 	jal	sin.2516
"10101011110111100000000000000010",	-- 9655: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 9656: 	lw	%ra, [%sp + 1]
"10010011110000010000000000000000",	-- 9657: 	lf	%f1, [%sp + 0]
"10110000000111100000000000000001",	-- 9658: 	sf	%f0, [%sp + 1]
"00001100001000000000000000000000",	-- 9659: 	movf	%f0, %f1
"00111111111111100000000000000010",	-- 9660: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9661: 	addi	%sp, %sp, 3
"01011000000000000000010010011000",	-- 9662: 	jal	cos.2518
"10101011110111100000000000000011",	-- 9663: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9664: 	lw	%ra, [%sp + 2]
"10010011110000010000000000000001",	-- 9665: 	lf	%f1, [%sp + 1]
"11101100001000000000000000000000",	-- 9666: 	divf	%f0, %f1, %f0
"01001111111000000000000000000000",	-- 9667: 	jr	%ra
	-- adjust_position.3000:
"11101000000000000000000000000000",	-- 9668: 	mulf	%f0, %f0, %f0
"00010100000000101100110011001101",	-- 9669: 	llif	%f2, 0.100000
"00010000000000100011110111001100",	-- 9670: 	lhif	%f2, 0.100000
"11100000000000100000000000000000",	-- 9671: 	addf	%f0, %f0, %f2
"10110000001111100000000000000000",	-- 9672: 	sf	%f1, [%sp + 0]
"00111111111111100000000000000001",	-- 9673: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 9674: 	addi	%sp, %sp, 2
"01011000000000000010101000110000",	-- 9675: 	jal	yj_sqrt
"10101011110111100000000000000010",	-- 9676: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 9677: 	lw	%ra, [%sp + 1]
"00010100000000010000000000000000",	-- 9678: 	llif	%f1, 1.000000
"00010000000000010011111110000000",	-- 9679: 	lhif	%f1, 1.000000
"11101100001000000000100000000000",	-- 9680: 	divf	%f1, %f1, %f0
"10110000000111100000000000000001",	-- 9681: 	sf	%f0, [%sp + 1]
"00001100001000000000000000000000",	-- 9682: 	movf	%f0, %f1
"00111111111111100000000000000010",	-- 9683: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9684: 	addi	%sp, %sp, 3
"01011000000000000000010010011110",	-- 9685: 	jal	atan.2520
"10101011110111100000000000000011",	-- 9686: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9687: 	lw	%ra, [%sp + 2]
"10010011110000010000000000000000",	-- 9688: 	lf	%f1, [%sp + 0]
"11101000000000010000000000000000",	-- 9689: 	mulf	%f0, %f0, %f1
"00111111111111100000000000000010",	-- 9690: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 9691: 	addi	%sp, %sp, 3
"01011000000000000010010110110011",	-- 9692: 	jal	tan.2998
"10101011110111100000000000000011",	-- 9693: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 9694: 	lw	%ra, [%sp + 2]
"10010011110000010000000000000001",	-- 9695: 	lf	%f1, [%sp + 1]
"11101000000000010000000000000000",	-- 9696: 	mulf	%f0, %f0, %f1
"01001111111000000000000000000000",	-- 9697: 	jr	%ra
	-- calc_dirvec.3003:
"00111011011001000000000000000001",	-- 9698: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000101",	-- 9699: 	lli	%r5, 5
"00110000101000010000000011011111",	-- 9700: 	bgt	%r5, %r1, bgt_else.9266
"00111100011111100000000000000000",	-- 9701: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 9702: 	sw	%r2, [%sp + 1]
"00111100100111100000000000000010",	-- 9703: 	sw	%r4, [%sp + 2]
"10110000000111100000000000000011",	-- 9704: 	sf	%f0, [%sp + 3]
"10110000001111100000000000000100",	-- 9705: 	sf	%f1, [%sp + 4]
"00111111111111100000000000000101",	-- 9706: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 9707: 	addi	%sp, %sp, 6
"01011000000000000000010011110001",	-- 9708: 	jal	fsqr.2530
"10101011110111100000000000000110",	-- 9709: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 9710: 	lw	%ra, [%sp + 5]
"10010011110000010000000000000100",	-- 9711: 	lf	%f1, [%sp + 4]
"10110000000111100000000000000101",	-- 9712: 	sf	%f0, [%sp + 5]
"00001100001000000000000000000000",	-- 9713: 	movf	%f0, %f1
"00111111111111100000000000000110",	-- 9714: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 9715: 	addi	%sp, %sp, 7
"01011000000000000000010011110001",	-- 9716: 	jal	fsqr.2530
"10101011110111100000000000000111",	-- 9717: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 9718: 	lw	%ra, [%sp + 6]
"10010011110000010000000000000101",	-- 9719: 	lf	%f1, [%sp + 5]
"11100000001000000000000000000000",	-- 9720: 	addf	%f0, %f1, %f0
"00010100000000010000000000000000",	-- 9721: 	llif	%f1, 1.000000
"00010000000000010011111110000000",	-- 9722: 	lhif	%f1, 1.000000
"11100000000000010000000000000000",	-- 9723: 	addf	%f0, %f0, %f1
"00111111111111100000000000000110",	-- 9724: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 9725: 	addi	%sp, %sp, 7
"01011000000000000010101000110000",	-- 9726: 	jal	yj_sqrt
"10101011110111100000000000000111",	-- 9727: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 9728: 	lw	%ra, [%sp + 6]
"10010011110000010000000000000011",	-- 9729: 	lf	%f1, [%sp + 3]
"11101100001000000000100000000000",	-- 9730: 	divf	%f1, %f1, %f0
"10010011110000100000000000000100",	-- 9731: 	lf	%f2, [%sp + 4]
"11101100010000000001000000000000",	-- 9732: 	divf	%f2, %f2, %f0
"00010100000000110000000000000000",	-- 9733: 	llif	%f3, 1.000000
"00010000000000110011111110000000",	-- 9734: 	lhif	%f3, 1.000000
"11101100011000000000000000000000",	-- 9735: 	divf	%f0, %f3, %f0
"00111011110000010000000000000001",	-- 9736: 	lw	%r1, [%sp + 1]
"00111011110000100000000000000010",	-- 9737: 	lw	%r2, [%sp + 2]
"10000100010000010000100000000000",	-- 9738: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 9739: 	lw	%r1, [%r1 + 0]
"00111011110000100000000000000000",	-- 9740: 	lw	%r2, [%sp + 0]
"10000100001000100001100000000000",	-- 9741: 	add	%r3, %r1, %r2
"00111000011000110000000000000000",	-- 9742: 	lw	%r3, [%r3 + 0]
"00111100001111100000000000000110",	-- 9743: 	sw	%r1, [%sp + 6]
"10110000000111100000000000000111",	-- 9744: 	sf	%f0, [%sp + 7]
"10110000010111100000000000001000",	-- 9745: 	sf	%f2, [%sp + 8]
"10110000001111100000000000001001",	-- 9746: 	sf	%f1, [%sp + 9]
"10000100000000110000100000000000",	-- 9747: 	add	%r1, %r0, %r3
"00111111111111100000000000001010",	-- 9748: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 9749: 	addi	%sp, %sp, 11
"01011000000000000000011010111100",	-- 9750: 	jal	d_vec.2683
"10101011110111100000000000001011",	-- 9751: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 9752: 	lw	%ra, [%sp + 10]
"10010011110000000000000000001001",	-- 9753: 	lf	%f0, [%sp + 9]
"10010011110000010000000000001000",	-- 9754: 	lf	%f1, [%sp + 8]
"10010011110000100000000000000111",	-- 9755: 	lf	%f2, [%sp + 7]
"00111111111111100000000000001010",	-- 9756: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 9757: 	addi	%sp, %sp, 11
"01011000000000000000010100100110",	-- 9758: 	jal	vecset.2576
"10101011110111100000000000001011",	-- 9759: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 9760: 	lw	%ra, [%sp + 10]
"11001100000000010000000000101000",	-- 9761: 	lli	%r1, 40
"00111011110000100000000000000000",	-- 9762: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 9763: 	add	%r1, %r2, %r1
"00111011110000110000000000000110",	-- 9764: 	lw	%r3, [%sp + 6]
"10000100011000010000100000000000",	-- 9765: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 9766: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001010",	-- 9767: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 9768: 	addi	%sp, %sp, 11
"01011000000000000000011010111100",	-- 9769: 	jal	d_vec.2683
"10101011110111100000000000001011",	-- 9770: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 9771: 	lw	%ra, [%sp + 10]
"10010011110000000000000000001000",	-- 9772: 	lf	%f0, [%sp + 8]
"00111100001111100000000000001010",	-- 9773: 	sw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 9774: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 9775: 	addi	%sp, %sp, 12
"01011000000000000010101001010001",	-- 9776: 	jal	yj_fneg
"10101011110111100000000000001100",	-- 9777: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9778: 	lw	%ra, [%sp + 11]
"00001100000000100000000000000000",	-- 9779: 	movf	%f2, %f0
"10010011110000000000000000001001",	-- 9780: 	lf	%f0, [%sp + 9]
"10010011110000010000000000000111",	-- 9781: 	lf	%f1, [%sp + 7]
"00111011110000010000000000001010",	-- 9782: 	lw	%r1, [%sp + 10]
"00111111111111100000000000001011",	-- 9783: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 9784: 	addi	%sp, %sp, 12
"01011000000000000000010100100110",	-- 9785: 	jal	vecset.2576
"10101011110111100000000000001100",	-- 9786: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9787: 	lw	%ra, [%sp + 11]
"11001100000000010000000001010000",	-- 9788: 	lli	%r1, 80
"00111011110000100000000000000000",	-- 9789: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 9790: 	add	%r1, %r2, %r1
"00111011110000110000000000000110",	-- 9791: 	lw	%r3, [%sp + 6]
"10000100011000010000100000000000",	-- 9792: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 9793: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001011",	-- 9794: 	sw	%ra, [%sp + 11]
"10100111110111100000000000001100",	-- 9795: 	addi	%sp, %sp, 12
"01011000000000000000011010111100",	-- 9796: 	jal	d_vec.2683
"10101011110111100000000000001100",	-- 9797: 	subi	%sp, %sp, 12
"00111011110111110000000000001011",	-- 9798: 	lw	%ra, [%sp + 11]
"10010011110000000000000000001001",	-- 9799: 	lf	%f0, [%sp + 9]
"00111100001111100000000000001011",	-- 9800: 	sw	%r1, [%sp + 11]
"00111111111111100000000000001100",	-- 9801: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 9802: 	addi	%sp, %sp, 13
"01011000000000000010101001010001",	-- 9803: 	jal	yj_fneg
"10101011110111100000000000001101",	-- 9804: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 9805: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001000",	-- 9806: 	lf	%f1, [%sp + 8]
"10110000000111100000000000001100",	-- 9807: 	sf	%f0, [%sp + 12]
"00001100001000000000000000000000",	-- 9808: 	movf	%f0, %f1
"00111111111111100000000000001101",	-- 9809: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 9810: 	addi	%sp, %sp, 14
"01011000000000000010101001010001",	-- 9811: 	jal	yj_fneg
"10101011110111100000000000001110",	-- 9812: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 9813: 	lw	%ra, [%sp + 13]
"00001100000000100000000000000000",	-- 9814: 	movf	%f2, %f0
"10010011110000000000000000000111",	-- 9815: 	lf	%f0, [%sp + 7]
"10010011110000010000000000001100",	-- 9816: 	lf	%f1, [%sp + 12]
"00111011110000010000000000001011",	-- 9817: 	lw	%r1, [%sp + 11]
"00111111111111100000000000001101",	-- 9818: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 9819: 	addi	%sp, %sp, 14
"01011000000000000000010100100110",	-- 9820: 	jal	vecset.2576
"10101011110111100000000000001110",	-- 9821: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 9822: 	lw	%ra, [%sp + 13]
"11001100000000010000000000000001",	-- 9823: 	lli	%r1, 1
"00111011110000100000000000000000",	-- 9824: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 9825: 	add	%r1, %r2, %r1
"00111011110000110000000000000110",	-- 9826: 	lw	%r3, [%sp + 6]
"10000100011000010000100000000000",	-- 9827: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 9828: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000001101",	-- 9829: 	sw	%ra, [%sp + 13]
"10100111110111100000000000001110",	-- 9830: 	addi	%sp, %sp, 14
"01011000000000000000011010111100",	-- 9831: 	jal	d_vec.2683
"10101011110111100000000000001110",	-- 9832: 	subi	%sp, %sp, 14
"00111011110111110000000000001101",	-- 9833: 	lw	%ra, [%sp + 13]
"10010011110000000000000000001001",	-- 9834: 	lf	%f0, [%sp + 9]
"00111100001111100000000000001101",	-- 9835: 	sw	%r1, [%sp + 13]
"00111111111111100000000000001110",	-- 9836: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 9837: 	addi	%sp, %sp, 15
"01011000000000000010101001010001",	-- 9838: 	jal	yj_fneg
"10101011110111100000000000001111",	-- 9839: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 9840: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001000",	-- 9841: 	lf	%f1, [%sp + 8]
"10110000000111100000000000001110",	-- 9842: 	sf	%f0, [%sp + 14]
"00001100001000000000000000000000",	-- 9843: 	movf	%f0, %f1
"00111111111111100000000000001111",	-- 9844: 	sw	%ra, [%sp + 15]
"10100111110111100000000000010000",	-- 9845: 	addi	%sp, %sp, 16
"01011000000000000010101001010001",	-- 9846: 	jal	yj_fneg
"10101011110111100000000000010000",	-- 9847: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 9848: 	lw	%ra, [%sp + 15]
"10010011110000010000000000000111",	-- 9849: 	lf	%f1, [%sp + 7]
"10110000000111100000000000001111",	-- 9850: 	sf	%f0, [%sp + 15]
"00001100001000000000000000000000",	-- 9851: 	movf	%f0, %f1
"00111111111111100000000000010000",	-- 9852: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 9853: 	addi	%sp, %sp, 17
"01011000000000000010101001010001",	-- 9854: 	jal	yj_fneg
"10101011110111100000000000010001",	-- 9855: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 9856: 	lw	%ra, [%sp + 16]
"00001100000000100000000000000000",	-- 9857: 	movf	%f2, %f0
"10010011110000000000000000001110",	-- 9858: 	lf	%f0, [%sp + 14]
"10010011110000010000000000001111",	-- 9859: 	lf	%f1, [%sp + 15]
"00111011110000010000000000001101",	-- 9860: 	lw	%r1, [%sp + 13]
"00111111111111100000000000010000",	-- 9861: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 9862: 	addi	%sp, %sp, 17
"01011000000000000000010100100110",	-- 9863: 	jal	vecset.2576
"10101011110111100000000000010001",	-- 9864: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 9865: 	lw	%ra, [%sp + 16]
"11001100000000010000000000101001",	-- 9866: 	lli	%r1, 41
"00111011110000100000000000000000",	-- 9867: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 9868: 	add	%r1, %r2, %r1
"00111011110000110000000000000110",	-- 9869: 	lw	%r3, [%sp + 6]
"10000100011000010000100000000000",	-- 9870: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 9871: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000010000",	-- 9872: 	sw	%ra, [%sp + 16]
"10100111110111100000000000010001",	-- 9873: 	addi	%sp, %sp, 17
"01011000000000000000011010111100",	-- 9874: 	jal	d_vec.2683
"10101011110111100000000000010001",	-- 9875: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 9876: 	lw	%ra, [%sp + 16]
"10010011110000000000000000001001",	-- 9877: 	lf	%f0, [%sp + 9]
"00111100001111100000000000010000",	-- 9878: 	sw	%r1, [%sp + 16]
"00111111111111100000000000010001",	-- 9879: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 9880: 	addi	%sp, %sp, 18
"01011000000000000010101001010001",	-- 9881: 	jal	yj_fneg
"10101011110111100000000000010010",	-- 9882: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 9883: 	lw	%ra, [%sp + 17]
"10010011110000010000000000000111",	-- 9884: 	lf	%f1, [%sp + 7]
"10110000000111100000000000010001",	-- 9885: 	sf	%f0, [%sp + 17]
"00001100001000000000000000000000",	-- 9886: 	movf	%f0, %f1
"00111111111111100000000000010010",	-- 9887: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 9888: 	addi	%sp, %sp, 19
"01011000000000000010101001010001",	-- 9889: 	jal	yj_fneg
"10101011110111100000000000010011",	-- 9890: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 9891: 	lw	%ra, [%sp + 18]
"00001100000000010000000000000000",	-- 9892: 	movf	%f1, %f0
"10010011110000000000000000010001",	-- 9893: 	lf	%f0, [%sp + 17]
"10010011110000100000000000001000",	-- 9894: 	lf	%f2, [%sp + 8]
"00111011110000010000000000010000",	-- 9895: 	lw	%r1, [%sp + 16]
"00111111111111100000000000010010",	-- 9896: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 9897: 	addi	%sp, %sp, 19
"01011000000000000000010100100110",	-- 9898: 	jal	vecset.2576
"10101011110111100000000000010011",	-- 9899: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 9900: 	lw	%ra, [%sp + 18]
"11001100000000010000000001010001",	-- 9901: 	lli	%r1, 81
"00111011110000100000000000000000",	-- 9902: 	lw	%r2, [%sp + 0]
"10000100010000010000100000000000",	-- 9903: 	add	%r1, %r2, %r1
"00111011110000100000000000000110",	-- 9904: 	lw	%r2, [%sp + 6]
"10000100010000010000100000000000",	-- 9905: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 9906: 	lw	%r1, [%r1 + 0]
"00111111111111100000000000010010",	-- 9907: 	sw	%ra, [%sp + 18]
"10100111110111100000000000010011",	-- 9908: 	addi	%sp, %sp, 19
"01011000000000000000011010111100",	-- 9909: 	jal	d_vec.2683
"10101011110111100000000000010011",	-- 9910: 	subi	%sp, %sp, 19
"00111011110111110000000000010010",	-- 9911: 	lw	%ra, [%sp + 18]
"10010011110000000000000000000111",	-- 9912: 	lf	%f0, [%sp + 7]
"00111100001111100000000000010010",	-- 9913: 	sw	%r1, [%sp + 18]
"00111111111111100000000000010011",	-- 9914: 	sw	%ra, [%sp + 19]
"10100111110111100000000000010100",	-- 9915: 	addi	%sp, %sp, 20
"01011000000000000010101001010001",	-- 9916: 	jal	yj_fneg
"10101011110111100000000000010100",	-- 9917: 	subi	%sp, %sp, 20
"00111011110111110000000000010011",	-- 9918: 	lw	%ra, [%sp + 19]
"10010011110000010000000000001001",	-- 9919: 	lf	%f1, [%sp + 9]
"10010011110000100000000000001000",	-- 9920: 	lf	%f2, [%sp + 8]
"00111011110000010000000000010010",	-- 9921: 	lw	%r1, [%sp + 18]
"01010100000000000000010100100110",	-- 9922: 	j	vecset.2576
	-- bgt_else.9266:
"10110000010111100000000000010011",	-- 9923: 	sf	%f2, [%sp + 19]
"00111100011111100000000000000000",	-- 9924: 	sw	%r3, [%sp + 0]
"00111100010111100000000000000001",	-- 9925: 	sw	%r2, [%sp + 1]
"00111111011111100000000000010100",	-- 9926: 	sw	%r27, [%sp + 20]
"10110000011111100000000000010101",	-- 9927: 	sf	%f3, [%sp + 21]
"00111100001111100000000000010110",	-- 9928: 	sw	%r1, [%sp + 22]
"00001100001000000000000000000000",	-- 9929: 	movf	%f0, %f1
"00001100010000010000000000000000",	-- 9930: 	movf	%f1, %f2
"00111111111111100000000000010111",	-- 9931: 	sw	%ra, [%sp + 23]
"10100111110111100000000000011000",	-- 9932: 	addi	%sp, %sp, 24
"01011000000000000010010111000100",	-- 9933: 	jal	adjust_position.3000
"10101011110111100000000000011000",	-- 9934: 	subi	%sp, %sp, 24
"00111011110111110000000000010111",	-- 9935: 	lw	%ra, [%sp + 23]
"11001100000000010000000000000001",	-- 9936: 	lli	%r1, 1
"00111011110000100000000000010110",	-- 9937: 	lw	%r2, [%sp + 22]
"10000100010000010000100000000000",	-- 9938: 	add	%r1, %r2, %r1
"10010011110000010000000000010101",	-- 9939: 	lf	%f1, [%sp + 21]
"10110000000111100000000000010111",	-- 9940: 	sf	%f0, [%sp + 23]
"00111100001111100000000000011000",	-- 9941: 	sw	%r1, [%sp + 24]
"00111111111111100000000000011001",	-- 9942: 	sw	%ra, [%sp + 25]
"10100111110111100000000000011010",	-- 9943: 	addi	%sp, %sp, 26
"01011000000000000010010111000100",	-- 9944: 	jal	adjust_position.3000
"10101011110111100000000000011010",	-- 9945: 	subi	%sp, %sp, 26
"00111011110111110000000000011001",	-- 9946: 	lw	%ra, [%sp + 25]
"00001100000000010000000000000000",	-- 9947: 	movf	%f1, %f0
"10010011110000000000000000010111",	-- 9948: 	lf	%f0, [%sp + 23]
"10010011110000100000000000010011",	-- 9949: 	lf	%f2, [%sp + 19]
"10010011110000110000000000010101",	-- 9950: 	lf	%f3, [%sp + 21]
"00111011110000010000000000011000",	-- 9951: 	lw	%r1, [%sp + 24]
"00111011110000100000000000000001",	-- 9952: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000000",	-- 9953: 	lw	%r3, [%sp + 0]
"00111011110110110000000000010100",	-- 9954: 	lw	%r27, [%sp + 20]
"00111011011110100000000000000000",	-- 9955: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 9956: 	jr	%r26
	-- calc_dirvecs.3011:
"00111011011001000000000000000001",	-- 9957: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 9958: 	lli	%r5, 0
"00110000101000010000000001010011",	-- 9959: 	bgt	%r5, %r1, bgt_else.9267
"00111111011111100000000000000000",	-- 9960: 	sw	%r27, [%sp + 0]
"00111100001111100000000000000001",	-- 9961: 	sw	%r1, [%sp + 1]
"10110000000111100000000000000010",	-- 9962: 	sf	%f0, [%sp + 2]
"00111100011111100000000000000011",	-- 9963: 	sw	%r3, [%sp + 3]
"00111100010111100000000000000100",	-- 9964: 	sw	%r2, [%sp + 4]
"00111100100111100000000000000101",	-- 9965: 	sw	%r4, [%sp + 5]
"00111111111111100000000000000110",	-- 9966: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 9967: 	addi	%sp, %sp, 7
"01011000000000000010101000101100",	-- 9968: 	jal	yj_float_of_int
"10101011110111100000000000000111",	-- 9969: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 9970: 	lw	%ra, [%sp + 6]
"00010100000000011100110011001101",	-- 9971: 	llif	%f1, 0.200000
"00010000000000010011111001001100",	-- 9972: 	lhif	%f1, 0.200000
"11101000000000010000000000000000",	-- 9973: 	mulf	%f0, %f0, %f1
"00010100000000010110011001100110",	-- 9974: 	llif	%f1, 0.900000
"00010000000000010011111101100110",	-- 9975: 	lhif	%f1, 0.900000
"11100100000000010001000000000000",	-- 9976: 	subf	%f2, %f0, %f1
"11001100000000010000000000000000",	-- 9977: 	lli	%r1, 0
"00010100000000000000000000000000",	-- 9978: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 9979: 	lhif	%f0, 0.000000
"00010100000000010000000000000000",	-- 9980: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 9981: 	lhif	%f1, 0.000000
"10010011110000110000000000000010",	-- 9982: 	lf	%f3, [%sp + 2]
"00111011110000100000000000000100",	-- 9983: 	lw	%r2, [%sp + 4]
"00111011110000110000000000000011",	-- 9984: 	lw	%r3, [%sp + 3]
"00111011110110110000000000000101",	-- 9985: 	lw	%r27, [%sp + 5]
"00111111111111100000000000000110",	-- 9986: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 9987: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 9988: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 9989: 	jalr	%r26
"10101011110111100000000000000111",	-- 9990: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 9991: 	lw	%ra, [%sp + 6]
"00111011110000010000000000000001",	-- 9992: 	lw	%r1, [%sp + 1]
"00111111111111100000000000000110",	-- 9993: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 9994: 	addi	%sp, %sp, 7
"01011000000000000010101000101100",	-- 9995: 	jal	yj_float_of_int
"10101011110111100000000000000111",	-- 9996: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 9997: 	lw	%ra, [%sp + 6]
"00010100000000011100110011001101",	-- 9998: 	llif	%f1, 0.200000
"00010000000000010011111001001100",	-- 9999: 	lhif	%f1, 0.200000
"11101000000000010000000000000000",	-- 10000: 	mulf	%f0, %f0, %f1
"00010100000000011100110011001101",	-- 10001: 	llif	%f1, 0.100000
"00010000000000010011110111001100",	-- 10002: 	lhif	%f1, 0.100000
"11100000000000010001000000000000",	-- 10003: 	addf	%f2, %f0, %f1
"11001100000000010000000000000000",	-- 10004: 	lli	%r1, 0
"00010100000000000000000000000000",	-- 10005: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 10006: 	lhif	%f0, 0.000000
"00010100000000010000000000000000",	-- 10007: 	llif	%f1, 0.000000
"00010000000000010000000000000000",	-- 10008: 	lhif	%f1, 0.000000
"11001100000000100000000000000010",	-- 10009: 	lli	%r2, 2
"00111011110000110000000000000011",	-- 10010: 	lw	%r3, [%sp + 3]
"10000100011000100001000000000000",	-- 10011: 	add	%r2, %r3, %r2
"10010011110000110000000000000010",	-- 10012: 	lf	%f3, [%sp + 2]
"00111011110001000000000000000100",	-- 10013: 	lw	%r4, [%sp + 4]
"00111011110110110000000000000101",	-- 10014: 	lw	%r27, [%sp + 5]
"10000100000000100001100000000000",	-- 10015: 	add	%r3, %r0, %r2
"10000100000001000001000000000000",	-- 10016: 	add	%r2, %r0, %r4
"00111111111111100000000000000110",	-- 10017: 	sw	%ra, [%sp + 6]
"00111011011110100000000000000000",	-- 10018: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000111",	-- 10019: 	addi	%sp, %sp, 7
"01010011010000000000000000000000",	-- 10020: 	jalr	%r26
"10101011110111100000000000000111",	-- 10021: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 10022: 	lw	%ra, [%sp + 6]
"11001100000000010000000000000001",	-- 10023: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 10024: 	lw	%r2, [%sp + 1]
"10001000010000010000100000000000",	-- 10025: 	sub	%r1, %r2, %r1
"11001100000000100000000000000001",	-- 10026: 	lli	%r2, 1
"00111011110000110000000000000100",	-- 10027: 	lw	%r3, [%sp + 4]
"00111100001111100000000000000110",	-- 10028: 	sw	%r1, [%sp + 6]
"10000100000000110000100000000000",	-- 10029: 	add	%r1, %r0, %r3
"00111111111111100000000000000111",	-- 10030: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 10031: 	addi	%sp, %sp, 8
"01011000000000000000010100011111",	-- 10032: 	jal	add_mod5.2573
"10101011110111100000000000001000",	-- 10033: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 10034: 	lw	%ra, [%sp + 7]
"10000100000000010001000000000000",	-- 10035: 	add	%r2, %r0, %r1
"10010011110000000000000000000010",	-- 10036: 	lf	%f0, [%sp + 2]
"00111011110000010000000000000110",	-- 10037: 	lw	%r1, [%sp + 6]
"00111011110000110000000000000011",	-- 10038: 	lw	%r3, [%sp + 3]
"00111011110110110000000000000000",	-- 10039: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10040: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10041: 	jr	%r26
	-- bgt_else.9267:
"01001111111000000000000000000000",	-- 10042: 	jr	%ra
	-- calc_dirvec_rows.3016:
"00111011011001000000000000000001",	-- 10043: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 10044: 	lli	%r5, 0
"00110000101000010000000000101111",	-- 10045: 	bgt	%r5, %r1, bgt_else.9269
"00111111011111100000000000000000",	-- 10046: 	sw	%r27, [%sp + 0]
"00111100001111100000000000000001",	-- 10047: 	sw	%r1, [%sp + 1]
"00111100011111100000000000000010",	-- 10048: 	sw	%r3, [%sp + 2]
"00111100010111100000000000000011",	-- 10049: 	sw	%r2, [%sp + 3]
"00111100100111100000000000000100",	-- 10050: 	sw	%r4, [%sp + 4]
"00111111111111100000000000000101",	-- 10051: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 10052: 	addi	%sp, %sp, 6
"01011000000000000010101000101100",	-- 10053: 	jal	yj_float_of_int
"10101011110111100000000000000110",	-- 10054: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 10055: 	lw	%ra, [%sp + 5]
"00010100000000011100110011001101",	-- 10056: 	llif	%f1, 0.200000
"00010000000000010011111001001100",	-- 10057: 	lhif	%f1, 0.200000
"11101000000000010000000000000000",	-- 10058: 	mulf	%f0, %f0, %f1
"00010100000000010110011001100110",	-- 10059: 	llif	%f1, 0.900000
"00010000000000010011111101100110",	-- 10060: 	lhif	%f1, 0.900000
"11100100000000010000000000000000",	-- 10061: 	subf	%f0, %f0, %f1
"11001100000000010000000000000100",	-- 10062: 	lli	%r1, 4
"00111011110000100000000000000011",	-- 10063: 	lw	%r2, [%sp + 3]
"00111011110000110000000000000010",	-- 10064: 	lw	%r3, [%sp + 2]
"00111011110110110000000000000100",	-- 10065: 	lw	%r27, [%sp + 4]
"00111111111111100000000000000101",	-- 10066: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 10067: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 10068: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 10069: 	jalr	%r26
"10101011110111100000000000000110",	-- 10070: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 10071: 	lw	%ra, [%sp + 5]
"11001100000000010000000000000001",	-- 10072: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 10073: 	lw	%r2, [%sp + 1]
"10001000010000010000100000000000",	-- 10074: 	sub	%r1, %r2, %r1
"11001100000000100000000000000010",	-- 10075: 	lli	%r2, 2
"00111011110000110000000000000011",	-- 10076: 	lw	%r3, [%sp + 3]
"00111100001111100000000000000101",	-- 10077: 	sw	%r1, [%sp + 5]
"10000100000000110000100000000000",	-- 10078: 	add	%r1, %r0, %r3
"00111111111111100000000000000110",	-- 10079: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 10080: 	addi	%sp, %sp, 7
"01011000000000000000010100011111",	-- 10081: 	jal	add_mod5.2573
"10101011110111100000000000000111",	-- 10082: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 10083: 	lw	%ra, [%sp + 6]
"10000100000000010001000000000000",	-- 10084: 	add	%r2, %r0, %r1
"11001100000000010000000000000100",	-- 10085: 	lli	%r1, 4
"00111011110000110000000000000010",	-- 10086: 	lw	%r3, [%sp + 2]
"10000100011000010001100000000000",	-- 10087: 	add	%r3, %r3, %r1
"00111011110000010000000000000101",	-- 10088: 	lw	%r1, [%sp + 5]
"00111011110110110000000000000000",	-- 10089: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10090: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10091: 	jr	%r26
	-- bgt_else.9269:
"01001111111000000000000000000000",	-- 10092: 	jr	%ra
	-- create_dirvec.3020:
"00111011011000010000000000000001",	-- 10093: 	lw	%r1, [%r27 + 1]
"11001100000000100000000000000011",	-- 10094: 	lli	%r2, 3
"00010100000000000000000000000000",	-- 10095: 	llif	%f0, 0.000000
"00010000000000000000000000000000",	-- 10096: 	lhif	%f0, 0.000000
"00111100001111100000000000000000",	-- 10097: 	sw	%r1, [%sp + 0]
"10000100000000100000100000000000",	-- 10098: 	add	%r1, %r0, %r2
"00111111111111100000000000000001",	-- 10099: 	sw	%ra, [%sp + 1]
"10100111110111100000000000000010",	-- 10100: 	addi	%sp, %sp, 2
"01011000000000000010101000100100",	-- 10101: 	jal	yj_create_float_array
"10101011110111100000000000000010",	-- 10102: 	subi	%sp, %sp, 2
"00111011110111110000000000000001",	-- 10103: 	lw	%ra, [%sp + 1]
"10000100000000010001000000000000",	-- 10104: 	add	%r2, %r0, %r1
"11001100000000010000000000000000",	-- 10105: 	lli	%r1, 0
"00111011110000110000000000000000",	-- 10106: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 10107: 	add	%r1, %r3, %r1
"00111000001000010000000000000000",	-- 10108: 	lw	%r1, [%r1 + 0]
"00111100010111100000000000000001",	-- 10109: 	sw	%r2, [%sp + 1]
"00111111111111100000000000000010",	-- 10110: 	sw	%ra, [%sp + 2]
"10100111110111100000000000000011",	-- 10111: 	addi	%sp, %sp, 3
"01011000000000000010101000011100",	-- 10112: 	jal	yj_create_array
"10101011110111100000000000000011",	-- 10113: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 10114: 	lw	%ra, [%sp + 2]
"10000100000111010001000000000000",	-- 10115: 	add	%r2, %r0, %hp
"10100111101111010000000000000010",	-- 10116: 	addi	%hp, %hp, 2
"00111100001000100000000000000001",	-- 10117: 	sw	%r1, [%r2 + 1]
"00111011110000010000000000000001",	-- 10118: 	lw	%r1, [%sp + 1]
"00111100001000100000000000000000",	-- 10119: 	sw	%r1, [%r2 + 0]
"10000100000000100000100000000000",	-- 10120: 	add	%r1, %r0, %r2
"01001111111000000000000000000000",	-- 10121: 	jr	%ra
	-- create_dirvec_elements.3022:
"00111011011000110000000000000001",	-- 10122: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 10123: 	lli	%r4, 0
"00110000100000100000000000010101",	-- 10124: 	bgt	%r4, %r2, bgt_else.9271
"00111111011111100000000000000000",	-- 10125: 	sw	%r27, [%sp + 0]
"00111100010111100000000000000001",	-- 10126: 	sw	%r2, [%sp + 1]
"00111100001111100000000000000010",	-- 10127: 	sw	%r1, [%sp + 2]
"10000100000000111101100000000000",	-- 10128: 	add	%r27, %r0, %r3
"00111111111111100000000000000011",	-- 10129: 	sw	%ra, [%sp + 3]
"00111011011110100000000000000000",	-- 10130: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000100",	-- 10131: 	addi	%sp, %sp, 4
"01010011010000000000000000000000",	-- 10132: 	jalr	%r26
"10101011110111100000000000000100",	-- 10133: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 10134: 	lw	%ra, [%sp + 3]
"00111011110000100000000000000001",	-- 10135: 	lw	%r2, [%sp + 1]
"00111011110000110000000000000010",	-- 10136: 	lw	%r3, [%sp + 2]
"10000100011000100010000000000000",	-- 10137: 	add	%r4, %r3, %r2
"00111100001001000000000000000000",	-- 10138: 	sw	%r1, [%r4 + 0]
"11001100000000010000000000000001",	-- 10139: 	lli	%r1, 1
"10001000010000010001000000000000",	-- 10140: 	sub	%r2, %r2, %r1
"00111011110110110000000000000000",	-- 10141: 	lw	%r27, [%sp + 0]
"10000100000000110000100000000000",	-- 10142: 	add	%r1, %r0, %r3
"00111011011110100000000000000000",	-- 10143: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10144: 	jr	%r26
	-- bgt_else.9271:
"01001111111000000000000000000000",	-- 10145: 	jr	%ra
	-- create_dirvecs.3025:
"00111011011000100000000000000011",	-- 10146: 	lw	%r2, [%r27 + 3]
"00111011011000110000000000000010",	-- 10147: 	lw	%r3, [%r27 + 2]
"00111011011001000000000000000001",	-- 10148: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 10149: 	lli	%r5, 0
"00110000101000010000000000101010",	-- 10150: 	bgt	%r5, %r1, bgt_else.9273
"11001100000001010000000001111000",	-- 10151: 	lli	%r5, 120
"00111111011111100000000000000000",	-- 10152: 	sw	%r27, [%sp + 0]
"00111100011111100000000000000001",	-- 10153: 	sw	%r3, [%sp + 1]
"00111100001111100000000000000010",	-- 10154: 	sw	%r1, [%sp + 2]
"00111100010111100000000000000011",	-- 10155: 	sw	%r2, [%sp + 3]
"00111100101111100000000000000100",	-- 10156: 	sw	%r5, [%sp + 4]
"10000100000001001101100000000000",	-- 10157: 	add	%r27, %r0, %r4
"00111111111111100000000000000101",	-- 10158: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 10159: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 10160: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 10161: 	jalr	%r26
"10101011110111100000000000000110",	-- 10162: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 10163: 	lw	%ra, [%sp + 5]
"10000100000000010001000000000000",	-- 10164: 	add	%r2, %r0, %r1
"00111011110000010000000000000100",	-- 10165: 	lw	%r1, [%sp + 4]
"00111111111111100000000000000101",	-- 10166: 	sw	%ra, [%sp + 5]
"10100111110111100000000000000110",	-- 10167: 	addi	%sp, %sp, 6
"01011000000000000010101000011100",	-- 10168: 	jal	yj_create_array
"10101011110111100000000000000110",	-- 10169: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 10170: 	lw	%ra, [%sp + 5]
"00111011110000100000000000000010",	-- 10171: 	lw	%r2, [%sp + 2]
"00111011110000110000000000000011",	-- 10172: 	lw	%r3, [%sp + 3]
"10000100011000100010000000000000",	-- 10173: 	add	%r4, %r3, %r2
"00111100001001000000000000000000",	-- 10174: 	sw	%r1, [%r4 + 0]
"10000100011000100000100000000000",	-- 10175: 	add	%r1, %r3, %r2
"00111000001000010000000000000000",	-- 10176: 	lw	%r1, [%r1 + 0]
"11001100000000110000000001110110",	-- 10177: 	lli	%r3, 118
"00111011110110110000000000000001",	-- 10178: 	lw	%r27, [%sp + 1]
"10000100000000110001000000000000",	-- 10179: 	add	%r2, %r0, %r3
"00111111111111100000000000000101",	-- 10180: 	sw	%ra, [%sp + 5]
"00111011011110100000000000000000",	-- 10181: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000110",	-- 10182: 	addi	%sp, %sp, 6
"01010011010000000000000000000000",	-- 10183: 	jalr	%r26
"10101011110111100000000000000110",	-- 10184: 	subi	%sp, %sp, 6
"00111011110111110000000000000101",	-- 10185: 	lw	%ra, [%sp + 5]
"11001100000000010000000000000001",	-- 10186: 	lli	%r1, 1
"00111011110000100000000000000010",	-- 10187: 	lw	%r2, [%sp + 2]
"10001000010000010000100000000000",	-- 10188: 	sub	%r1, %r2, %r1
"00111011110110110000000000000000",	-- 10189: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10190: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10191: 	jr	%r26
	-- bgt_else.9273:
"01001111111000000000000000000000",	-- 10192: 	jr	%ra
	-- init_dirvec_constants.3027:
"00111011011000110000000000000001",	-- 10193: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 10194: 	lli	%r4, 0
"00110000100000100000000000010101",	-- 10195: 	bgt	%r4, %r2, bgt_else.9275
"10000100001000100010000000000000",	-- 10196: 	add	%r4, %r1, %r2
"00111000100001000000000000000000",	-- 10197: 	lw	%r4, [%r4 + 0]
"00111100001111100000000000000000",	-- 10198: 	sw	%r1, [%sp + 0]
"00111111011111100000000000000001",	-- 10199: 	sw	%r27, [%sp + 1]
"00111100010111100000000000000010",	-- 10200: 	sw	%r2, [%sp + 2]
"10000100000001000000100000000000",	-- 10201: 	add	%r1, %r0, %r4
"10000100000000111101100000000000",	-- 10202: 	add	%r27, %r0, %r3
"00111111111111100000000000000011",	-- 10203: 	sw	%ra, [%sp + 3]
"00111011011110100000000000000000",	-- 10204: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000100",	-- 10205: 	addi	%sp, %sp, 4
"01010011010000000000000000000000",	-- 10206: 	jalr	%r26
"10101011110111100000000000000100",	-- 10207: 	subi	%sp, %sp, 4
"00111011110111110000000000000011",	-- 10208: 	lw	%ra, [%sp + 3]
"11001100000000010000000000000001",	-- 10209: 	lli	%r1, 1
"00111011110000100000000000000010",	-- 10210: 	lw	%r2, [%sp + 2]
"10001000010000010001000000000000",	-- 10211: 	sub	%r2, %r2, %r1
"00111011110000010000000000000000",	-- 10212: 	lw	%r1, [%sp + 0]
"00111011110110110000000000000001",	-- 10213: 	lw	%r27, [%sp + 1]
"00111011011110100000000000000000",	-- 10214: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10215: 	jr	%r26
	-- bgt_else.9275:
"01001111111000000000000000000000",	-- 10216: 	jr	%ra
	-- init_vecset_constants.3030:
"00111011011000100000000000000010",	-- 10217: 	lw	%r2, [%r27 + 2]
"00111011011000110000000000000001",	-- 10218: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000000",	-- 10219: 	lli	%r4, 0
"00110000100000010000000000010101",	-- 10220: 	bgt	%r4, %r1, bgt_else.9277
"10000100011000010001100000000000",	-- 10221: 	add	%r3, %r3, %r1
"00111000011000110000000000000000",	-- 10222: 	lw	%r3, [%r3 + 0]
"11001100000001000000000001110111",	-- 10223: 	lli	%r4, 119
"00111111011111100000000000000000",	-- 10224: 	sw	%r27, [%sp + 0]
"00111100001111100000000000000001",	-- 10225: 	sw	%r1, [%sp + 1]
"10000100000000110000100000000000",	-- 10226: 	add	%r1, %r0, %r3
"10000100000000101101100000000000",	-- 10227: 	add	%r27, %r0, %r2
"10000100000001000001000000000000",	-- 10228: 	add	%r2, %r0, %r4
"00111111111111100000000000000010",	-- 10229: 	sw	%ra, [%sp + 2]
"00111011011110100000000000000000",	-- 10230: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000011",	-- 10231: 	addi	%sp, %sp, 3
"01010011010000000000000000000000",	-- 10232: 	jalr	%r26
"10101011110111100000000000000011",	-- 10233: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 10234: 	lw	%ra, [%sp + 2]
"11001100000000010000000000000001",	-- 10235: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 10236: 	lw	%r2, [%sp + 1]
"10001000010000010000100000000000",	-- 10237: 	sub	%r1, %r2, %r1
"00111011110110110000000000000000",	-- 10238: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10239: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10240: 	jr	%r26
	-- bgt_else.9277:
"01001111111000000000000000000000",	-- 10241: 	jr	%ra
	-- init_dirvecs.3032:
"00111011011000010000000000000011",	-- 10242: 	lw	%r1, [%r27 + 3]
"00111011011000100000000000000010",	-- 10243: 	lw	%r2, [%r27 + 2]
"00111011011000110000000000000001",	-- 10244: 	lw	%r3, [%r27 + 1]
"11001100000001000000000000000100",	-- 10245: 	lli	%r4, 4
"00111100001111100000000000000000",	-- 10246: 	sw	%r1, [%sp + 0]
"00111100011111100000000000000001",	-- 10247: 	sw	%r3, [%sp + 1]
"10000100000001000000100000000000",	-- 10248: 	add	%r1, %r0, %r4
"10000100000000101101100000000000",	-- 10249: 	add	%r27, %r0, %r2
"00111111111111100000000000000010",	-- 10250: 	sw	%ra, [%sp + 2]
"00111011011110100000000000000000",	-- 10251: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000011",	-- 10252: 	addi	%sp, %sp, 3
"01010011010000000000000000000000",	-- 10253: 	jalr	%r26
"10101011110111100000000000000011",	-- 10254: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 10255: 	lw	%ra, [%sp + 2]
"11001100000000010000000000001001",	-- 10256: 	lli	%r1, 9
"11001100000000100000000000000000",	-- 10257: 	lli	%r2, 0
"11001100000000110000000000000000",	-- 10258: 	lli	%r3, 0
"00111011110110110000000000000001",	-- 10259: 	lw	%r27, [%sp + 1]
"00111111111111100000000000000010",	-- 10260: 	sw	%ra, [%sp + 2]
"00111011011110100000000000000000",	-- 10261: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000000011",	-- 10262: 	addi	%sp, %sp, 3
"01010011010000000000000000000000",	-- 10263: 	jalr	%r26
"10101011110111100000000000000011",	-- 10264: 	subi	%sp, %sp, 3
"00111011110111110000000000000010",	-- 10265: 	lw	%ra, [%sp + 2]
"11001100000000010000000000000100",	-- 10266: 	lli	%r1, 4
"00111011110110110000000000000000",	-- 10267: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10268: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10269: 	jr	%r26
	-- add_reflection.3034:
"00111011011000110000000000000011",	-- 10270: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 10271: 	lw	%r4, [%r27 + 2]
"00111011011110110000000000000001",	-- 10272: 	lw	%r27, [%r27 + 1]
"00111100001111100000000000000000",	-- 10273: 	sw	%r1, [%sp + 0]
"00111100100111100000000000000001",	-- 10274: 	sw	%r4, [%sp + 1]
"00111100010111100000000000000010",	-- 10275: 	sw	%r2, [%sp + 2]
"10110000000111100000000000000011",	-- 10276: 	sf	%f0, [%sp + 3]
"00111100011111100000000000000100",	-- 10277: 	sw	%r3, [%sp + 4]
"10110000011111100000000000000101",	-- 10278: 	sf	%f3, [%sp + 5]
"10110000010111100000000000000110",	-- 10279: 	sf	%f2, [%sp + 6]
"10110000001111100000000000000111",	-- 10280: 	sf	%f1, [%sp + 7]
"00111111111111100000000000001000",	-- 10281: 	sw	%ra, [%sp + 8]
"00111011011110100000000000000000",	-- 10282: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001001",	-- 10283: 	addi	%sp, %sp, 9
"01010011010000000000000000000000",	-- 10284: 	jalr	%r26
"10101011110111100000000000001001",	-- 10285: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 10286: 	lw	%ra, [%sp + 8]
"00111100001111100000000000001000",	-- 10287: 	sw	%r1, [%sp + 8]
"00111111111111100000000000001001",	-- 10288: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 10289: 	addi	%sp, %sp, 10
"01011000000000000000011010111100",	-- 10290: 	jal	d_vec.2683
"10101011110111100000000000001010",	-- 10291: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 10292: 	lw	%ra, [%sp + 9]
"10010011110000000000000000000111",	-- 10293: 	lf	%f0, [%sp + 7]
"10010011110000010000000000000110",	-- 10294: 	lf	%f1, [%sp + 6]
"10010011110000100000000000000101",	-- 10295: 	lf	%f2, [%sp + 5]
"00111111111111100000000000001001",	-- 10296: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 10297: 	addi	%sp, %sp, 10
"01011000000000000000010100100110",	-- 10298: 	jal	vecset.2576
"10101011110111100000000000001010",	-- 10299: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 10300: 	lw	%ra, [%sp + 9]
"00111011110000010000000000001000",	-- 10301: 	lw	%r1, [%sp + 8]
"00111011110110110000000000000100",	-- 10302: 	lw	%r27, [%sp + 4]
"00111111111111100000000000001001",	-- 10303: 	sw	%ra, [%sp + 9]
"00111011011110100000000000000000",	-- 10304: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001010",	-- 10305: 	addi	%sp, %sp, 10
"01010011010000000000000000000000",	-- 10306: 	jalr	%r26
"10101011110111100000000000001010",	-- 10307: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 10308: 	lw	%ra, [%sp + 9]
"10000100000111010000100000000000",	-- 10309: 	add	%r1, %r0, %hp
"10100111101111010000000000000011",	-- 10310: 	addi	%hp, %hp, 3
"10010011110000000000000000000011",	-- 10311: 	lf	%f0, [%sp + 3]
"10110000000000010000000000000010",	-- 10312: 	sf	%f0, [%r1 + 2]
"00111011110000100000000000001000",	-- 10313: 	lw	%r2, [%sp + 8]
"00111100010000010000000000000001",	-- 10314: 	sw	%r2, [%r1 + 1]
"00111011110000100000000000000010",	-- 10315: 	lw	%r2, [%sp + 2]
"00111100010000010000000000000000",	-- 10316: 	sw	%r2, [%r1 + 0]
"00111011110000100000000000000000",	-- 10317: 	lw	%r2, [%sp + 0]
"00111011110000110000000000000001",	-- 10318: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 10319: 	add	%r2, %r3, %r2
"00111100001000100000000000000000",	-- 10320: 	sw	%r1, [%r2 + 0]
"01001111111000000000000000000000",	-- 10321: 	jr	%ra
	-- setup_rect_reflection.3041:
"00111011011000110000000000000011",	-- 10322: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 10323: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 10324: 	lw	%r5, [%r27 + 1]
"11001100000001100000000000000100",	-- 10325: 	lli	%r6, 4
"10001100001001100000100000000000",	-- 10326: 	mul	%r1, %r1, %r6
"11001100000001100000000000000000",	-- 10327: 	lli	%r6, 0
"10000100011001100011000000000000",	-- 10328: 	add	%r6, %r3, %r6
"00111000110001100000000000000000",	-- 10329: 	lw	%r6, [%r6 + 0]
"00010100000000000000000000000000",	-- 10330: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 10331: 	lhif	%f0, 1.000000
"00111100011111100000000000000000",	-- 10332: 	sw	%r3, [%sp + 0]
"00111100110111100000000000000001",	-- 10333: 	sw	%r6, [%sp + 1]
"00111100101111100000000000000010",	-- 10334: 	sw	%r5, [%sp + 2]
"00111100001111100000000000000011",	-- 10335: 	sw	%r1, [%sp + 3]
"00111100100111100000000000000100",	-- 10336: 	sw	%r4, [%sp + 4]
"10110000000111100000000000000101",	-- 10337: 	sf	%f0, [%sp + 5]
"10000100000000100000100000000000",	-- 10338: 	add	%r1, %r0, %r2
"00111111111111100000000000000110",	-- 10339: 	sw	%ra, [%sp + 6]
"10100111110111100000000000000111",	-- 10340: 	addi	%sp, %sp, 7
"01011000000000000000011001111010",	-- 10341: 	jal	o_diffuse.2646
"10101011110111100000000000000111",	-- 10342: 	subi	%sp, %sp, 7
"00111011110111110000000000000110",	-- 10343: 	lw	%ra, [%sp + 6]
"10010011110000010000000000000101",	-- 10344: 	lf	%f1, [%sp + 5]
"11100100001000000000000000000000",	-- 10345: 	subf	%f0, %f1, %f0
"11001100000000010000000000000000",	-- 10346: 	lli	%r1, 0
"00111011110000100000000000000100",	-- 10347: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 10348: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 10349: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000110",	-- 10350: 	sf	%f0, [%sp + 6]
"00001100001000000000000000000000",	-- 10351: 	movf	%f0, %f1
"00111111111111100000000000000111",	-- 10352: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 10353: 	addi	%sp, %sp, 8
"01011000000000000010101001010001",	-- 10354: 	jal	yj_fneg
"10101011110111100000000000001000",	-- 10355: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 10356: 	lw	%ra, [%sp + 7]
"11001100000000010000000000000001",	-- 10357: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 10358: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 10359: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 10360: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000000111",	-- 10361: 	sf	%f0, [%sp + 7]
"00001100001000000000000000000000",	-- 10362: 	movf	%f0, %f1
"00111111111111100000000000001000",	-- 10363: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 10364: 	addi	%sp, %sp, 9
"01011000000000000010101001010001",	-- 10365: 	jal	yj_fneg
"10101011110111100000000000001001",	-- 10366: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 10367: 	lw	%ra, [%sp + 8]
"11001100000000010000000000000010",	-- 10368: 	lli	%r1, 2
"00111011110000100000000000000100",	-- 10369: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 10370: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 10371: 	lf	%f1, [%r1 + 0]
"10110000000111100000000000001000",	-- 10372: 	sf	%f0, [%sp + 8]
"00001100001000000000000000000000",	-- 10373: 	movf	%f0, %f1
"00111111111111100000000000001001",	-- 10374: 	sw	%ra, [%sp + 9]
"10100111110111100000000000001010",	-- 10375: 	addi	%sp, %sp, 10
"01011000000000000010101001010001",	-- 10376: 	jal	yj_fneg
"10101011110111100000000000001010",	-- 10377: 	subi	%sp, %sp, 10
"00111011110111110000000000001001",	-- 10378: 	lw	%ra, [%sp + 9]
"00001100000000110000000000000000",	-- 10379: 	movf	%f3, %f0
"11001100000000010000000000000001",	-- 10380: 	lli	%r1, 1
"00111011110000100000000000000011",	-- 10381: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 10382: 	add	%r1, %r2, %r1
"11001100000000110000000000000000",	-- 10383: 	lli	%r3, 0
"00111011110001000000000000000100",	-- 10384: 	lw	%r4, [%sp + 4]
"10000100100000110001100000000000",	-- 10385: 	add	%r3, %r4, %r3
"10010000011000010000000000000000",	-- 10386: 	lf	%f1, [%r3 + 0]
"10010011110000000000000000000110",	-- 10387: 	lf	%f0, [%sp + 6]
"10010011110000100000000000001000",	-- 10388: 	lf	%f2, [%sp + 8]
"00111011110000110000000000000001",	-- 10389: 	lw	%r3, [%sp + 1]
"00111011110110110000000000000010",	-- 10390: 	lw	%r27, [%sp + 2]
"10110000011111100000000000001001",	-- 10391: 	sf	%f3, [%sp + 9]
"10000100000000010001000000000000",	-- 10392: 	add	%r2, %r0, %r1
"10000100000000110000100000000000",	-- 10393: 	add	%r1, %r0, %r3
"00111111111111100000000000001010",	-- 10394: 	sw	%ra, [%sp + 10]
"00111011011110100000000000000000",	-- 10395: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001011",	-- 10396: 	addi	%sp, %sp, 11
"01010011010000000000000000000000",	-- 10397: 	jalr	%r26
"10101011110111100000000000001011",	-- 10398: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 10399: 	lw	%ra, [%sp + 10]
"11001100000000010000000000000001",	-- 10400: 	lli	%r1, 1
"00111011110000100000000000000001",	-- 10401: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 10402: 	add	%r1, %r2, %r1
"11001100000000110000000000000010",	-- 10403: 	lli	%r3, 2
"00111011110001000000000000000011",	-- 10404: 	lw	%r4, [%sp + 3]
"10000100100000110001100000000000",	-- 10405: 	add	%r3, %r4, %r3
"11001100000001010000000000000001",	-- 10406: 	lli	%r5, 1
"00111011110001100000000000000100",	-- 10407: 	lw	%r6, [%sp + 4]
"10000100110001010010100000000000",	-- 10408: 	add	%r5, %r6, %r5
"10010000101000100000000000000000",	-- 10409: 	lf	%f2, [%r5 + 0]
"10010011110000000000000000000110",	-- 10410: 	lf	%f0, [%sp + 6]
"10010011110000010000000000000111",	-- 10411: 	lf	%f1, [%sp + 7]
"10010011110000110000000000001001",	-- 10412: 	lf	%f3, [%sp + 9]
"00111011110110110000000000000010",	-- 10413: 	lw	%r27, [%sp + 2]
"10000100000000110001000000000000",	-- 10414: 	add	%r2, %r0, %r3
"00111111111111100000000000001010",	-- 10415: 	sw	%ra, [%sp + 10]
"00111011011110100000000000000000",	-- 10416: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001011",	-- 10417: 	addi	%sp, %sp, 11
"01010011010000000000000000000000",	-- 10418: 	jalr	%r26
"10101011110111100000000000001011",	-- 10419: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 10420: 	lw	%ra, [%sp + 10]
"11001100000000010000000000000010",	-- 10421: 	lli	%r1, 2
"00111011110000100000000000000001",	-- 10422: 	lw	%r2, [%sp + 1]
"10000100010000010000100000000000",	-- 10423: 	add	%r1, %r2, %r1
"11001100000000110000000000000011",	-- 10424: 	lli	%r3, 3
"00111011110001000000000000000011",	-- 10425: 	lw	%r4, [%sp + 3]
"10000100100000110001100000000000",	-- 10426: 	add	%r3, %r4, %r3
"11001100000001000000000000000010",	-- 10427: 	lli	%r4, 2
"00111011110001010000000000000100",	-- 10428: 	lw	%r5, [%sp + 4]
"10000100101001000010000000000000",	-- 10429: 	add	%r4, %r5, %r4
"10010000100000110000000000000000",	-- 10430: 	lf	%f3, [%r4 + 0]
"10010011110000000000000000000110",	-- 10431: 	lf	%f0, [%sp + 6]
"10010011110000010000000000000111",	-- 10432: 	lf	%f1, [%sp + 7]
"10010011110000100000000000001000",	-- 10433: 	lf	%f2, [%sp + 8]
"00111011110110110000000000000010",	-- 10434: 	lw	%r27, [%sp + 2]
"10000100000000110001000000000000",	-- 10435: 	add	%r2, %r0, %r3
"00111111111111100000000000001010",	-- 10436: 	sw	%ra, [%sp + 10]
"00111011011110100000000000000000",	-- 10437: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001011",	-- 10438: 	addi	%sp, %sp, 11
"01010011010000000000000000000000",	-- 10439: 	jalr	%r26
"10101011110111100000000000001011",	-- 10440: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 10441: 	lw	%ra, [%sp + 10]
"11001100000000010000000000000000",	-- 10442: 	lli	%r1, 0
"11001100000000100000000000000011",	-- 10443: 	lli	%r2, 3
"00111011110000110000000000000001",	-- 10444: 	lw	%r3, [%sp + 1]
"10000100011000100001000000000000",	-- 10445: 	add	%r2, %r3, %r2
"00111011110000110000000000000000",	-- 10446: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 10447: 	add	%r1, %r3, %r1
"00111100010000010000000000000000",	-- 10448: 	sw	%r2, [%r1 + 0]
"01001111111000000000000000000000",	-- 10449: 	jr	%ra
	-- setup_surface_reflection.3044:
"00111011011000110000000000000011",	-- 10450: 	lw	%r3, [%r27 + 3]
"00111011011001000000000000000010",	-- 10451: 	lw	%r4, [%r27 + 2]
"00111011011001010000000000000001",	-- 10452: 	lw	%r5, [%r27 + 1]
"11001100000001100000000000000100",	-- 10453: 	lli	%r6, 4
"10001100001001100000100000000000",	-- 10454: 	mul	%r1, %r1, %r6
"11001100000001100000000000000001",	-- 10455: 	lli	%r6, 1
"10000100001001100000100000000000",	-- 10456: 	add	%r1, %r1, %r6
"11001100000001100000000000000000",	-- 10457: 	lli	%r6, 0
"10000100011001100011000000000000",	-- 10458: 	add	%r6, %r3, %r6
"00111000110001100000000000000000",	-- 10459: 	lw	%r6, [%r6 + 0]
"00010100000000000000000000000000",	-- 10460: 	llif	%f0, 1.000000
"00010000000000000011111110000000",	-- 10461: 	lhif	%f0, 1.000000
"00111100011111100000000000000000",	-- 10462: 	sw	%r3, [%sp + 0]
"00111100001111100000000000000001",	-- 10463: 	sw	%r1, [%sp + 1]
"00111100110111100000000000000010",	-- 10464: 	sw	%r6, [%sp + 2]
"00111100101111100000000000000011",	-- 10465: 	sw	%r5, [%sp + 3]
"00111100100111100000000000000100",	-- 10466: 	sw	%r4, [%sp + 4]
"00111100010111100000000000000101",	-- 10467: 	sw	%r2, [%sp + 5]
"10110000000111100000000000000110",	-- 10468: 	sf	%f0, [%sp + 6]
"10000100000000100000100000000000",	-- 10469: 	add	%r1, %r0, %r2
"00111111111111100000000000000111",	-- 10470: 	sw	%ra, [%sp + 7]
"10100111110111100000000000001000",	-- 10471: 	addi	%sp, %sp, 8
"01011000000000000000011001111010",	-- 10472: 	jal	o_diffuse.2646
"10101011110111100000000000001000",	-- 10473: 	subi	%sp, %sp, 8
"00111011110111110000000000000111",	-- 10474: 	lw	%ra, [%sp + 7]
"10010011110000010000000000000110",	-- 10475: 	lf	%f1, [%sp + 6]
"11100100001000000000000000000000",	-- 10476: 	subf	%f0, %f1, %f0
"00111011110000010000000000000101",	-- 10477: 	lw	%r1, [%sp + 5]
"10110000000111100000000000000111",	-- 10478: 	sf	%f0, [%sp + 7]
"00111111111111100000000000001000",	-- 10479: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 10480: 	addi	%sp, %sp, 9
"01011000000000000000011001101001",	-- 10481: 	jal	o_param_abc.2638
"10101011110111100000000000001001",	-- 10482: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 10483: 	lw	%ra, [%sp + 8]
"10000100000000010001000000000000",	-- 10484: 	add	%r2, %r0, %r1
"00111011110000010000000000000100",	-- 10485: 	lw	%r1, [%sp + 4]
"00111111111111100000000000001000",	-- 10486: 	sw	%ra, [%sp + 8]
"10100111110111100000000000001001",	-- 10487: 	addi	%sp, %sp, 9
"01011000000000000000010110100111",	-- 10488: 	jal	veciprod.2597
"10101011110111100000000000001001",	-- 10489: 	subi	%sp, %sp, 9
"00111011110111110000000000001000",	-- 10490: 	lw	%ra, [%sp + 8]
"00010100000000010000000000000000",	-- 10491: 	llif	%f1, 2.000000
"00010000000000010100000000000000",	-- 10492: 	lhif	%f1, 2.000000
"00111011110000010000000000000101",	-- 10493: 	lw	%r1, [%sp + 5]
"10110000000111100000000000001000",	-- 10494: 	sf	%f0, [%sp + 8]
"10110000001111100000000000001001",	-- 10495: 	sf	%f1, [%sp + 9]
"00111111111111100000000000001010",	-- 10496: 	sw	%ra, [%sp + 10]
"10100111110111100000000000001011",	-- 10497: 	addi	%sp, %sp, 11
"01011000000000000000011001011010",	-- 10498: 	jal	o_param_a.2632
"10101011110111100000000000001011",	-- 10499: 	subi	%sp, %sp, 11
"00111011110111110000000000001010",	-- 10500: 	lw	%ra, [%sp + 10]
"10010011110000010000000000001001",	-- 10501: 	lf	%f1, [%sp + 9]
"11101000001000000000000000000000",	-- 10502: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001000",	-- 10503: 	lf	%f1, [%sp + 8]
"11101000000000010000000000000000",	-- 10504: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000000",	-- 10505: 	lli	%r1, 0
"00111011110000100000000000000100",	-- 10506: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 10507: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 10508: 	lf	%f2, [%r1 + 0]
"11100100000000100000000000000000",	-- 10509: 	subf	%f0, %f0, %f2
"00010100000000100000000000000000",	-- 10510: 	llif	%f2, 2.000000
"00010000000000100100000000000000",	-- 10511: 	lhif	%f2, 2.000000
"00111011110000010000000000000101",	-- 10512: 	lw	%r1, [%sp + 5]
"10110000000111100000000000001010",	-- 10513: 	sf	%f0, [%sp + 10]
"10110000010111100000000000001011",	-- 10514: 	sf	%f2, [%sp + 11]
"00111111111111100000000000001100",	-- 10515: 	sw	%ra, [%sp + 12]
"10100111110111100000000000001101",	-- 10516: 	addi	%sp, %sp, 13
"01011000000000000000011001011111",	-- 10517: 	jal	o_param_b.2634
"10101011110111100000000000001101",	-- 10518: 	subi	%sp, %sp, 13
"00111011110111110000000000001100",	-- 10519: 	lw	%ra, [%sp + 12]
"10010011110000010000000000001011",	-- 10520: 	lf	%f1, [%sp + 11]
"11101000001000000000000000000000",	-- 10521: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001000",	-- 10522: 	lf	%f1, [%sp + 8]
"11101000000000010000000000000000",	-- 10523: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000001",	-- 10524: 	lli	%r1, 1
"00111011110000100000000000000100",	-- 10525: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 10526: 	add	%r1, %r2, %r1
"10010000001000100000000000000000",	-- 10527: 	lf	%f2, [%r1 + 0]
"11100100000000100000000000000000",	-- 10528: 	subf	%f0, %f0, %f2
"00010100000000100000000000000000",	-- 10529: 	llif	%f2, 2.000000
"00010000000000100100000000000000",	-- 10530: 	lhif	%f2, 2.000000
"00111011110000010000000000000101",	-- 10531: 	lw	%r1, [%sp + 5]
"10110000000111100000000000001100",	-- 10532: 	sf	%f0, [%sp + 12]
"10110000010111100000000000001101",	-- 10533: 	sf	%f2, [%sp + 13]
"00111111111111100000000000001110",	-- 10534: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 10535: 	addi	%sp, %sp, 15
"01011000000000000000011001100100",	-- 10536: 	jal	o_param_c.2636
"10101011110111100000000000001111",	-- 10537: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 10538: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001101",	-- 10539: 	lf	%f1, [%sp + 13]
"11101000001000000000000000000000",	-- 10540: 	mulf	%f0, %f1, %f0
"10010011110000010000000000001000",	-- 10541: 	lf	%f1, [%sp + 8]
"11101000000000010000000000000000",	-- 10542: 	mulf	%f0, %f0, %f1
"11001100000000010000000000000010",	-- 10543: 	lli	%r1, 2
"00111011110000100000000000000100",	-- 10544: 	lw	%r2, [%sp + 4]
"10000100010000010000100000000000",	-- 10545: 	add	%r1, %r2, %r1
"10010000001000010000000000000000",	-- 10546: 	lf	%f1, [%r1 + 0]
"11100100000000010001100000000000",	-- 10547: 	subf	%f3, %f0, %f1
"10010011110000000000000000000111",	-- 10548: 	lf	%f0, [%sp + 7]
"10010011110000010000000000001010",	-- 10549: 	lf	%f1, [%sp + 10]
"10010011110000100000000000001100",	-- 10550: 	lf	%f2, [%sp + 12]
"00111011110000010000000000000010",	-- 10551: 	lw	%r1, [%sp + 2]
"00111011110000100000000000000001",	-- 10552: 	lw	%r2, [%sp + 1]
"00111011110110110000000000000011",	-- 10553: 	lw	%r27, [%sp + 3]
"00111111111111100000000000001110",	-- 10554: 	sw	%ra, [%sp + 14]
"00111011011110100000000000000000",	-- 10555: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001111",	-- 10556: 	addi	%sp, %sp, 15
"01010011010000000000000000000000",	-- 10557: 	jalr	%r26
"10101011110111100000000000001111",	-- 10558: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 10559: 	lw	%ra, [%sp + 14]
"11001100000000010000000000000000",	-- 10560: 	lli	%r1, 0
"11001100000000100000000000000001",	-- 10561: 	lli	%r2, 1
"00111011110000110000000000000010",	-- 10562: 	lw	%r3, [%sp + 2]
"10000100011000100001000000000000",	-- 10563: 	add	%r2, %r3, %r2
"00111011110000110000000000000000",	-- 10564: 	lw	%r3, [%sp + 0]
"10000100011000010000100000000000",	-- 10565: 	add	%r1, %r3, %r1
"00111100010000010000000000000000",	-- 10566: 	sw	%r2, [%r1 + 0]
"01001111111000000000000000000000",	-- 10567: 	jr	%ra
	-- setup_reflections.3047:
"00111011011000100000000000000011",	-- 10568: 	lw	%r2, [%r27 + 3]
"00111011011000110000000000000010",	-- 10569: 	lw	%r3, [%r27 + 2]
"00111011011001000000000000000001",	-- 10570: 	lw	%r4, [%r27 + 1]
"11001100000001010000000000000000",	-- 10571: 	lli	%r5, 0
"00110000101000010000000000110101",	-- 10572: 	bgt	%r5, %r1, bgt_else.9282
"10000100100000010010000000000000",	-- 10573: 	add	%r4, %r4, %r1
"00111000100001000000000000000000",	-- 10574: 	lw	%r4, [%r4 + 0]
"00111100010111100000000000000000",	-- 10575: 	sw	%r2, [%sp + 0]
"00111100001111100000000000000001",	-- 10576: 	sw	%r1, [%sp + 1]
"00111100011111100000000000000010",	-- 10577: 	sw	%r3, [%sp + 2]
"00111100100111100000000000000011",	-- 10578: 	sw	%r4, [%sp + 3]
"10000100000001000000100000000000",	-- 10579: 	add	%r1, %r0, %r4
"00111111111111100000000000000100",	-- 10580: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 10581: 	addi	%sp, %sp, 5
"01011000000000000000011001010100",	-- 10582: 	jal	o_reflectiontype.2626
"10101011110111100000000000000101",	-- 10583: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 10584: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000010",	-- 10585: 	lli	%r2, 2
"00101000001000100000000000100110",	-- 10586: 	bneq	%r1, %r2, bneq_else.9283
"00111011110000010000000000000011",	-- 10587: 	lw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 10588: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 10589: 	addi	%sp, %sp, 5
"01011000000000000000011001111010",	-- 10590: 	jal	o_diffuse.2646
"10101011110111100000000000000101",	-- 10591: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 10592: 	lw	%ra, [%sp + 4]
"00010100000000010000000000000000",	-- 10593: 	llif	%f1, 1.000000
"00010000000000010011111110000000",	-- 10594: 	lhif	%f1, 1.000000
"00111111111111100000000000000100",	-- 10595: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 10596: 	addi	%sp, %sp, 5
"01011000000000000000010011110011",	-- 10597: 	jal	fless.2532
"10101011110111100000000000000101",	-- 10598: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 10599: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000000",	-- 10600: 	lli	%r2, 0
"00101000001000100000000000000010",	-- 10601: 	bneq	%r1, %r2, bneq_else.9284
"01001111111000000000000000000000",	-- 10602: 	jr	%ra
	-- bneq_else.9284:
"00111011110000010000000000000011",	-- 10603: 	lw	%r1, [%sp + 3]
"00111111111111100000000000000100",	-- 10604: 	sw	%ra, [%sp + 4]
"10100111110111100000000000000101",	-- 10605: 	addi	%sp, %sp, 5
"01011000000000000000011001010010",	-- 10606: 	jal	o_form.2624
"10101011110111100000000000000101",	-- 10607: 	subi	%sp, %sp, 5
"00111011110111110000000000000100",	-- 10608: 	lw	%ra, [%sp + 4]
"11001100000000100000000000000001",	-- 10609: 	lli	%r2, 1
"00101000001000100000000000000110",	-- 10610: 	bneq	%r1, %r2, bneq_else.9286
"00111011110000010000000000000001",	-- 10611: 	lw	%r1, [%sp + 1]
"00111011110000100000000000000011",	-- 10612: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000010",	-- 10613: 	lw	%r27, [%sp + 2]
"00111011011110100000000000000000",	-- 10614: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10615: 	jr	%r26
	-- bneq_else.9286:
"11001100000000100000000000000010",	-- 10616: 	lli	%r2, 2
"00101000001000100000000000000110",	-- 10617: 	bneq	%r1, %r2, bneq_else.9287
"00111011110000010000000000000001",	-- 10618: 	lw	%r1, [%sp + 1]
"00111011110000100000000000000011",	-- 10619: 	lw	%r2, [%sp + 3]
"00111011110110110000000000000000",	-- 10620: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10621: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10622: 	jr	%r26
	-- bneq_else.9287:
"01001111111000000000000000000000",	-- 10623: 	jr	%ra
	-- bneq_else.9283:
"01001111111000000000000000000000",	-- 10624: 	jr	%ra
	-- bgt_else.9282:
"01001111111000000000000000000000",	-- 10625: 	jr	%ra
	-- rt.3049:
"00111011011000110000000000001110",	-- 10626: 	lw	%r3, [%r27 + 14]
"00111011011001000000000000001101",	-- 10627: 	lw	%r4, [%r27 + 13]
"00111011011001010000000000001100",	-- 10628: 	lw	%r5, [%r27 + 12]
"00111011011001100000000000001011",	-- 10629: 	lw	%r6, [%r27 + 11]
"00111011011001110000000000001010",	-- 10630: 	lw	%r7, [%r27 + 10]
"00111011011010000000000000001001",	-- 10631: 	lw	%r8, [%r27 + 9]
"00111011011010010000000000001000",	-- 10632: 	lw	%r9, [%r27 + 8]
"00111011011010100000000000000111",	-- 10633: 	lw	%r10, [%r27 + 7]
"00111011011010110000000000000110",	-- 10634: 	lw	%r11, [%r27 + 6]
"00111011011011000000000000000101",	-- 10635: 	lw	%r12, [%r27 + 5]
"00111011011011010000000000000100",	-- 10636: 	lw	%r13, [%r27 + 4]
"00111011011011100000000000000011",	-- 10637: 	lw	%r14, [%r27 + 3]
"00111011011011110000000000000010",	-- 10638: 	lw	%r15, [%r27 + 2]
"00111011011100000000000000000001",	-- 10639: 	lw	%r16, [%r27 + 1]
"11001100000100010000000000000000",	-- 10640: 	lli	%r17, 0
"10000101110100011000100000000000",	-- 10641: 	add	%r17, %r14, %r17
"00111100001100010000000000000000",	-- 10642: 	sw	%r1, [%r17 + 0]
"11001100000100010000000000000001",	-- 10643: 	lli	%r17, 1
"10000101110100010111000000000000",	-- 10644: 	add	%r14, %r14, %r17
"00111100010011100000000000000000",	-- 10645: 	sw	%r2, [%r14 + 0]
"11001100000011100000000000000000",	-- 10646: 	lli	%r14, 0
"01000000001100010000000000000001",	-- 10647: 	sra	%r17, %r1, 1
"10000101111011100111000000000000",	-- 10648: 	add	%r14, %r15, %r14
"00111110001011100000000000000000",	-- 10649: 	sw	%r17, [%r14 + 0]
"11001100000011100000000000000001",	-- 10650: 	lli	%r14, 1
"01000000010000100000000000000001",	-- 10651: 	sra	%r2, %r2, 1
"10000101111011100111000000000000",	-- 10652: 	add	%r14, %r15, %r14
"00111100010011100000000000000000",	-- 10653: 	sw	%r2, [%r14 + 0]
"11001100000000100000000000000000",	-- 10654: 	lli	%r2, 0
"00010100000000000000000000000000",	-- 10655: 	llif	%f0, 128.000000
"00010000000000000100001100000000",	-- 10656: 	lhif	%f0, 128.000000
"00111100111111100000000000000000",	-- 10657: 	sw	%r7, [%sp + 0]
"00111101001111100000000000000001",	-- 10658: 	sw	%r9, [%sp + 1]
"00111100100111100000000000000010",	-- 10659: 	sw	%r4, [%sp + 2]
"00111101010111100000000000000011",	-- 10660: 	sw	%r10, [%sp + 3]
"00111100101111100000000000000100",	-- 10661: 	sw	%r5, [%sp + 4]
"00111101100111100000000000000101",	-- 10662: 	sw	%r12, [%sp + 5]
"00111101011111100000000000000110",	-- 10663: 	sw	%r11, [%sp + 6]
"00111101101111100000000000000111",	-- 10664: 	sw	%r13, [%sp + 7]
"00111100011111100000000000001000",	-- 10665: 	sw	%r3, [%sp + 8]
"00111101000111100000000000001001",	-- 10666: 	sw	%r8, [%sp + 9]
"00111110000111100000000000001010",	-- 10667: 	sw	%r16, [%sp + 10]
"00111100010111100000000000001011",	-- 10668: 	sw	%r2, [%sp + 11]
"00111100110111100000000000001100",	-- 10669: 	sw	%r6, [%sp + 12]
"10110000000111100000000000001101",	-- 10670: 	sf	%f0, [%sp + 13]
"00111111111111100000000000001110",	-- 10671: 	sw	%ra, [%sp + 14]
"10100111110111100000000000001111",	-- 10672: 	addi	%sp, %sp, 15
"01011000000000000010101000101100",	-- 10673: 	jal	yj_float_of_int
"10101011110111100000000000001111",	-- 10674: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 10675: 	lw	%ra, [%sp + 14]
"10010011110000010000000000001101",	-- 10676: 	lf	%f1, [%sp + 13]
"11101100001000000000000000000000",	-- 10677: 	divf	%f0, %f1, %f0
"00111011110000010000000000001011",	-- 10678: 	lw	%r1, [%sp + 11]
"00111011110000100000000000001100",	-- 10679: 	lw	%r2, [%sp + 12]
"10000100010000010000100000000000",	-- 10680: 	add	%r1, %r2, %r1
"10110000000000010000000000000000",	-- 10681: 	sf	%f0, [%r1 + 0]
"00111011110110110000000000001010",	-- 10682: 	lw	%r27, [%sp + 10]
"00111111111111100000000000001110",	-- 10683: 	sw	%ra, [%sp + 14]
"00111011011110100000000000000000",	-- 10684: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000001111",	-- 10685: 	addi	%sp, %sp, 15
"01010011010000000000000000000000",	-- 10686: 	jalr	%r26
"10101011110111100000000000001111",	-- 10687: 	subi	%sp, %sp, 15
"00111011110111110000000000001110",	-- 10688: 	lw	%ra, [%sp + 14]
"00111011110110110000000000001010",	-- 10689: 	lw	%r27, [%sp + 10]
"00111100001111100000000000001110",	-- 10690: 	sw	%r1, [%sp + 14]
"00111111111111100000000000001111",	-- 10691: 	sw	%ra, [%sp + 15]
"00111011011110100000000000000000",	-- 10692: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010000",	-- 10693: 	addi	%sp, %sp, 16
"01010011010000000000000000000000",	-- 10694: 	jalr	%r26
"10101011110111100000000000010000",	-- 10695: 	subi	%sp, %sp, 16
"00111011110111110000000000001111",	-- 10696: 	lw	%ra, [%sp + 15]
"00111011110110110000000000001010",	-- 10697: 	lw	%r27, [%sp + 10]
"00111100001111100000000000001111",	-- 10698: 	sw	%r1, [%sp + 15]
"00111111111111100000000000010000",	-- 10699: 	sw	%ra, [%sp + 16]
"00111011011110100000000000000000",	-- 10700: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010001",	-- 10701: 	addi	%sp, %sp, 17
"01010011010000000000000000000000",	-- 10702: 	jalr	%r26
"10101011110111100000000000010001",	-- 10703: 	subi	%sp, %sp, 17
"00111011110111110000000000010000",	-- 10704: 	lw	%ra, [%sp + 16]
"00111011110110110000000000001001",	-- 10705: 	lw	%r27, [%sp + 9]
"00111100001111100000000000010000",	-- 10706: 	sw	%r1, [%sp + 16]
"00111111111111100000000000010001",	-- 10707: 	sw	%ra, [%sp + 17]
"00111011011110100000000000000000",	-- 10708: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010010",	-- 10709: 	addi	%sp, %sp, 18
"01010011010000000000000000000000",	-- 10710: 	jalr	%r26
"10101011110111100000000000010010",	-- 10711: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10712: 	lw	%ra, [%sp + 17]
"00111011110110110000000000001000",	-- 10713: 	lw	%r27, [%sp + 8]
"00111111111111100000000000010001",	-- 10714: 	sw	%ra, [%sp + 17]
"00111011011110100000000000000000",	-- 10715: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010010",	-- 10716: 	addi	%sp, %sp, 18
"01010011010000000000000000000000",	-- 10717: 	jalr	%r26
"10101011110111100000000000010010",	-- 10718: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10719: 	lw	%ra, [%sp + 17]
"00111011110110110000000000000111",	-- 10720: 	lw	%r27, [%sp + 7]
"00111111111111100000000000010001",	-- 10721: 	sw	%ra, [%sp + 17]
"00111011011110100000000000000000",	-- 10722: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010010",	-- 10723: 	addi	%sp, %sp, 18
"01010011010000000000000000000000",	-- 10724: 	jalr	%r26
"10101011110111100000000000010010",	-- 10725: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10726: 	lw	%ra, [%sp + 17]
"00111011110000010000000000000110",	-- 10727: 	lw	%r1, [%sp + 6]
"00111111111111100000000000010001",	-- 10728: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 10729: 	addi	%sp, %sp, 18
"01011000000000000000011010111100",	-- 10730: 	jal	d_vec.2683
"10101011110111100000000000010010",	-- 10731: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10732: 	lw	%ra, [%sp + 17]
"00111011110000100000000000000101",	-- 10733: 	lw	%r2, [%sp + 5]
"00111111111111100000000000010001",	-- 10734: 	sw	%ra, [%sp + 17]
"10100111110111100000000000010010",	-- 10735: 	addi	%sp, %sp, 18
"01011000000000000000010100111101",	-- 10736: 	jal	veccpy.2586
"10101011110111100000000000010010",	-- 10737: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10738: 	lw	%ra, [%sp + 17]
"00111011110000010000000000000110",	-- 10739: 	lw	%r1, [%sp + 6]
"00111011110110110000000000000100",	-- 10740: 	lw	%r27, [%sp + 4]
"00111111111111100000000000010001",	-- 10741: 	sw	%ra, [%sp + 17]
"00111011011110100000000000000000",	-- 10742: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010010",	-- 10743: 	addi	%sp, %sp, 18
"01010011010000000000000000000000",	-- 10744: 	jalr	%r26
"10101011110111100000000000010010",	-- 10745: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10746: 	lw	%ra, [%sp + 17]
"11001100000000010000000000000000",	-- 10747: 	lli	%r1, 0
"00111011110000100000000000000011",	-- 10748: 	lw	%r2, [%sp + 3]
"10000100010000010000100000000000",	-- 10749: 	add	%r1, %r2, %r1
"00111000001000010000000000000000",	-- 10750: 	lw	%r1, [%r1 + 0]
"11001100000000100000000000000001",	-- 10751: 	lli	%r2, 1
"10001000001000100000100000000000",	-- 10752: 	sub	%r1, %r1, %r2
"00111011110110110000000000000010",	-- 10753: 	lw	%r27, [%sp + 2]
"00111111111111100000000000010001",	-- 10754: 	sw	%ra, [%sp + 17]
"00111011011110100000000000000000",	-- 10755: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010010",	-- 10756: 	addi	%sp, %sp, 18
"01010011010000000000000000000000",	-- 10757: 	jalr	%r26
"10101011110111100000000000010010",	-- 10758: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10759: 	lw	%ra, [%sp + 17]
"11001100000000100000000000000000",	-- 10760: 	lli	%r2, 0
"11001100000000110000000000000000",	-- 10761: 	lli	%r3, 0
"00111011110000010000000000001111",	-- 10762: 	lw	%r1, [%sp + 15]
"00111011110110110000000000000001",	-- 10763: 	lw	%r27, [%sp + 1]
"00111111111111100000000000010001",	-- 10764: 	sw	%ra, [%sp + 17]
"00111011011110100000000000000000",	-- 10765: 	lw	%r26, [%r27 + 0]
"10100111110111100000000000010010",	-- 10766: 	addi	%sp, %sp, 18
"01010011010000000000000000000000",	-- 10767: 	jalr	%r26
"10101011110111100000000000010010",	-- 10768: 	subi	%sp, %sp, 18
"00111011110111110000000000010001",	-- 10769: 	lw	%ra, [%sp + 17]
"11001100000000010000000000000000",	-- 10770: 	lli	%r1, 0
"11001100000001010000000000000010",	-- 10771: 	lli	%r5, 2
"00111011110000100000000000001110",	-- 10772: 	lw	%r2, [%sp + 14]
"00111011110000110000000000001111",	-- 10773: 	lw	%r3, [%sp + 15]
"00111011110001000000000000010000",	-- 10774: 	lw	%r4, [%sp + 16]
"00111011110110110000000000000000",	-- 10775: 	lw	%r27, [%sp + 0]
"00111011011110100000000000000000",	-- 10776: 	lw	%r26, [%r27 + 0]
"01001111010000000000000000000000",	-- 10777: 	jr	%r26
	-- yj_print_char:
"11010000001000000000000000000000",	-- 10778: 	sendc	%r1
"01001111111000000000000000000000",	-- 10779: 	jr	%ra
	-- yj_create_array:
"11001100000000110000000000000000",	-- 10780: 	lli	%r3, 0
	-- yj_create.loop:
"10000111101000110010000000000000",	-- 10781: 	add	%r4, %hp, %r3
"00111100010001000000000000000000",	-- 10782: 	sw	%r2, [%r4 + 0]
"10100100011000110000000000000001",	-- 10783: 	addi	%r3, %r3, 1
"00110000001000111111111111111101",	-- 10784: 	bgt	%r1, %r3, yj_create.loop
"10000100000111010000100000000000",	-- 10785: 	add	%r1, %r0, %hp
"10000111101000111110100000000000",	-- 10786: 	add	%hp, %hp, %r3
"01001111111000000000000000000000",	-- 10787: 	jr	%ra
	-- yj_create_float_array:
"11001100000000110000000000000000",	-- 10788: 	lli	%r3, 0
	-- yj_create_float.loop:
"10000111101000110010000000000000",	-- 10789: 	add	%r4, %hp, %r3
"10110000000001000000000000000000",	-- 10790: 	sf	%f0, [%r4 + 0]
"10100100011000110000000000000001",	-- 10791: 	addi	%r3, %r3, 1
"00110000001000111111111111111101",	-- 10792: 	bgt	%r1, %r3, yj_create_float.loop
"10000100000111010000100000000000",	-- 10793: 	add	%r1, %r0, %hp
"10000111101000111110100000000000",	-- 10794: 	add	%hp, %hp, %r3
"01001111111000000000000000000000",	-- 10795: 	jr	%ra
	-- yj_float_of_int:
"01100000001000000000000000000000",	-- 10796: 	itof	%f0, %r1
"01001111111000000000000000000000",	-- 10797: 	jr	%ra
	-- yj_int_of_float:
"01100100000000010000000000000000",	-- 10798: 	ftoi	%r1, %f0
"01001111111000000000000000000000",	-- 10799: 	jr	%ra
	-- yj_sqrt:
"11110000000000000000000000000000",	-- 10800: 	sqrt	%f0, %f0
"01001111111000000000000000000000",	-- 10801: 	jr	%ra
	-- yj_floor:
"11110100000000000000000000000000",	-- 10802: 	floor	%f0, %f0
"01001111111000000000000000000000",	-- 10803: 	jr	%ra
	-- yj_read_int:
"11001100000000010000000000000000",	-- 10804: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 10805: 	lli	%r2, 0
"11000100000000010000000000000000",	-- 10806: 	recv	%r1
"01001000001000010000000000001000",	-- 10807: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 10808: 	recv	%r2
"10011100001000100000100000000000",	-- 10809: 	xor	%r1, %r1, %r2
"01001000001000010000000000001000",	-- 10810: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 10811: 	recv	%r2
"10011100001000100000100000000000",	-- 10812: 	xor	%r1, %r1, %r2
"01001000001000010000000000001000",	-- 10813: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 10814: 	recv	%r2
"10011100001000100000100000000000",	-- 10815: 	xor	%r1, %r1, %r2
"01001111111000000000000000000000",	-- 10816: 	jr	%ra
	-- yj_read_float:
"11001100000000010000000000000000",	-- 10817: 	lli	%r1, 0
"11001100000000100000000000000000",	-- 10818: 	lli	%r2, 0
"11000100000000010000000000000000",	-- 10819: 	recv	%r1
"01001000001000010000000000001000",	-- 10820: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 10821: 	recv	%r2
"10011100001000100000100000000000",	-- 10822: 	xor	%r1, %r1, %r2
"01001000001000010000000000001000",	-- 10823: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 10824: 	recv	%r2
"10011100001000100000100000000000",	-- 10825: 	xor	%r1, %r1, %r2
"01001000001000010000000000001000",	-- 10826: 	sll	%r1, %r1, 8
"11000100000000100000000000000000",	-- 10827: 	recv	%r2
"10011100001000100000100000000000",	-- 10828: 	xor	%r1, %r1, %r2
"01111100001000000000000000000000",	-- 10829: 	movi2f	%f0, %r1
"01001111111000000000000000000000",	-- 10830: 	jr	%ra
	-- yj_fabs:
"11111000000000000000000000000000",	-- 10831: 	absf	%f0, %f0
"01001111111000000000000000000000",	-- 10832: 	jr	%ra
	-- yj_fneg:
"00011000000000000000000000000000",	-- 10833: 	negf	%f0, %f0
"01001111111000000000000000000000"	-- 10834: 	jr	%ra
);

signal shortened : std_logic_vector(6 downto 0):=(others=>'0');
begin  -- R_rom
  shortened<=addra(6 downto 0);
    douta<=rom(conv_integer(shortened));
end R_rom;
