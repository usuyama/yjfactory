library IEEE;
use IEEE.std_logic_1164.all;

library work;

package fdiv_table is

subtype vector is std_logic_vector(23 downto 0);
type vector2 is array (0 to 2047) of vector;
constant table : vector2 :=(
"111111111110000000000100",
"111111111100000000010000",
"111111111010000000100100",
"111111111000000001000000",
"111111110110000001100100",
"111111110100000010010000",
"111111110010000011000011",
"111111110000000011111111",
"111111101110000101000011",
"111111101100000110001110",
"111111101010000111100001",
"111111101000001000111101",
"111111100110001010100000",
"111111100100001100001011",
"111111100010001101111101",
"111111100000001111111000",
"111111011110010001111010",
"111111011100010100000101",
"111111011010010110010111",
"111111011000011000110001",
"111111010110011011010010",
"111111010100011101111011",
"111111010010100000101101",
"111111010000100011100101",
"111111001110100110100110",
"111111001100101001101110",
"111111001010101100111110",
"111111001000110000010110",
"111111000110110011110101",
"111111000100110111011100",
"111111000010111011001011",
"111111000000111111000001",
"111110111111000010111111",
"111110111101000111000100",
"111110111011001011010010",
"111110111001001111100110",
"111110110111010100000011",
"111110110101011000100111",
"111110110011011101010010",
"111110110001100010000101",
"111110101111100111000000",
"111110101101101100000010",
"111110101011110001001100",
"111110101001110110011101",
"111110100111111011110110",
"111110100110000001010110",
"111110100100000110111110",
"111110100010001100101101",
"111110100000010010100100",
"111110011110011000100010",
"111110011100011110100111",
"111110011010100100110100",
"111110011000101011001001",
"111110010110110001100100",
"111110010100111000001000",
"111110010010111110110010",
"111110010001000101100100",
"111110001111001100011101",
"111110001101010011011110",
"111110001011011010100110",
"111110001001100001110110",
"111110000111101001001100",
"111110000101110000101010",
"111110000011111000010000",
"111110000001111111111100",
"111110000000000111110000",
"111101111110001111101011",
"111101111100010111101110",
"111101111010011111110111",
"111101111000101000001000",
"111101110110110000100000",
"111101110100111001000000",
"111101110011000001100110",
"111101110001001010010100",
"111101101111010011001001",
"111101101101011100000101",
"111101101011100101001001",
"111101101001101110010011",
"111101100111110111100101",
"111101100110000000111110",
"111101100100001010011110",
"111101100010010100000101",
"111101100000011101110011",
"111101011110100111101000",
"111101011100110001100100",
"111101011010111011101000",
"111101011001000101110010",
"111101010111010000000100",
"111101010101011010011100",
"111101010011100100111100",
"111101010001101111100011",
"111101001111111010010001",
"111101001110000101000101",
"111101001100010000000001",
"111101001010011011000100",
"111101001000100110001101",
"111101000110110001011110",
"111101000100111100110110",
"111101000011001000010100",
"111101000001010011111010",
"111100111111011111100110",
"111100111101101011011010",
"111100111011110111010100",
"111100111010000011010101",
"111100111000001111011101",
"111100110110011011101100",
"111100110100101000000010",
"111100110010110100011111",
"111100110001000001000010",
"111100101111001101101101",
"111100101101011010011110",
"111100101011100111010110",
"111100101001110100010101",
"111100101000000001011011",
"111100100110001110100111",
"111100100100011011111011",
"111100100010101001010101",
"111100100000110110110110",
"111100011111000100011101",
"111100011101010010001100",
"111100011011100000000001",
"111100011001101101111101",
"111100010111111011111111",
"111100010110001010001001",
"111100010100011000011001",
"111100010010100110101111",
"111100010000110101001101",
"111100001111000011110001",
"111100001101010010011100",
"111100001011100001001101",
"111100001001110000000101",
"111100000111111111000100",
"111100000110001110001001",
"111100000100011101010101",
"111100000010101100101000",
"111100000000111100000001",
"111011111111001011100001",
"111011111101011011000111",
"111011111011101010110100",
"111011111001111010101000",
"111011111000001010100010",
"111011110110011010100010",
"111011110100101010101001",
"111011110010111010110111",
"111011110001001011001011",
"111011101111011011100110",
"111011101101101100000111",
"111011101011111100101111",
"111011101010001101011101",
"111011101000011110010010",
"111011100110101111001101",
"111011100101000000001111",
"111011100011010001010111",
"111011100001100010100110",
"111011011111110011111011",
"111011011110000101010110",
"111011011100010110111000",
"111011011010101000100000",
"111011011000111010001111",
"111011010111001100000100",
"111011010101011101111111",
"111011010011110000000001",
"111011010010000010001001",
"111011010000010100011000",
"111011001110100110101100",
"111011001100111001001000",
"111011001011001011101001",
"111011001001011110010001",
"111011000111110000111111",
"111011000110000011110100",
"111011000100010110101111",
"111011000010101001110000",
"111011000000111100110111",
"111010111111010000000101",
"111010111101100011011001",
"111010111011110110110011",
"111010111010001010010011",
"111010111000011101111010",
"111010110110110001100111",
"111010110101000101011010",
"111010110011011001010011",
"111010110001101101010010",
"111010110000000001011000",
"111010101110010101100100",
"111010101100101001110110",
"111010101010111110001110",
"111010101001010010101101",
"111010100111100111010001",
"111010100101111011111100",
"111010100100010000101101",
"111010100010100101100100",
"111010100000111010100001",
"111010011111001111100100",
"111010011101100100101101",
"111010011011111001111101",
"111010011010001111010010",
"111010011000100100101110",
"111010010110111010010000",
"111010010101001111110111",
"111010010011100101100101",
"111010010001111011011001",
"111010010000010001010011",
"111010001110100111010011",
"111010001100111101011001",
"111010001011010011100101",
"111010001001101001110111",
"111010001000000000001111",
"111010000110010110101100",
"111010000100101101010000",
"111010000011000011111010",
"111010000001011010101010",
"111001111111110001100000",
"111001111110001000011100",
"111001111100011111011110",
"111001111010110110100101",
"111001111001001101110011",
"111001110111100101000110",
"111001110101111100100000",
"111001110100010011111111",
"111001110010101011100100",
"111001110001000011010000",
"111001101111011011000001",
"111001101101110010111000",
"111001101100001010110100",
"111001101010100010110111",
"111001101000111010111111",
"111001100111010011001110",
"111001100101101011100010",
"111001100100000011111100",
"111001100010011100011100",
"111001100000110101000001",
"111001011111001101101101",
"111001011101100110011110",
"111001011011111111010101",
"111001011010011000010010",
"111001011000110001010100",
"111001010111001010011101",
"111001010101100011101011",
"111001010011111100111111",
"111001010010010110011000",
"111001010000101111111000",
"111001001111001001011101",
"111001001101100011000111",
"111001001011111100111000",
"111001001010010110101110",
"111001001000110000101010",
"111001000111001010101100",
"111001000101100100110011",
"111001000011111111000000",
"111001000010011001010010",
"111001000000110011101011",
"111000111111001110001001",
"111000111101101000101100",
"111000111100000011010110",
"111000111010011110000100",
"111000111000111000111001",
"111000110111010011110011",
"111000110101101110110011",
"111000110100001001111000",
"111000110010100101000011",
"111000110001000000010100",
"111000101111011011101010",
"111000101101110111000101",
"111000101100010010100111",
"111000101010101110001101",
"111000101001001001111010",
"111000100111100101101100",
"111000100110000001100011",
"111000100100011101100000",
"111000100010111001100011",
"111000100001010101101011",
"111000011111110001111000",
"111000011110001110001011",
"111000011100101010100100",
"111000011011000111000010",
"111000011001100011100101",
"111000011000000000001110",
"111000010110011100111101",
"111000010100111001110000",
"111000010011010110101010",
"111000010001110011101001",
"111000010000010000101101",
"111000001110101101110111",
"111000001101001011000110",
"111000001011101000011010",
"111000001010000101110100",
"111000001000100011010011",
"111000000111000000111000",
"111000000101011110100010",
"111000000011111100010010",
"111000000010011010000111",
"111000000000111000000001",
"110111111111010110000000",
"110111111101110100000101",
"110111111100010010010000",
"110111111010110000011111",
"110111111001001110110100",
"110111110111101101001111",
"110111110110001011101110",
"110111110100101010010011",
"110111110011001000111110",
"110111110001100111101101",
"110111110000000110100010",
"110111101110100101011100",
"110111101101000100011100",
"110111101011100011100000",
"110111101010000010101010",
"110111101000100001111010",
"110111100111000001001110",
"110111100101100000101000",
"110111100100000000000111",
"110111100010011111101011",
"110111100000111111010101",
"110111011111011111000011",
"110111011101111110110111",
"110111011100011110110000",
"110111011010111110101111",
"110111011001011110110010",
"110111010111111110111011",
"110111010110011111001001",
"110111010100111111011100",
"110111010011011111110100",
"110111010010000000010001",
"110111010000100000110100",
"110111001111000001011011",
"110111001101100010001000",
"110111001100000010111010",
"110111001010100011110001",
"110111001001000100101110",
"110111000111100101101111",
"110111000110000110110101",
"110111000100101000000001",
"110111000011001001010001",
"110111000001101010100111",
"110111000000001100000010",
"110110111110101101100010",
"110110111101001111000111",
"110110111011110000110001",
"110110111010010010100000",
"110110111000110100010100",
"110110110111010110001101",
"110110110101111000001100",
"110110110100011010001111",
"110110110010111100010111",
"110110110001011110100100",
"110110110000000000110111",
"110110101110100011001110",
"110110101101000101101010",
"110110101011101000001100",
"110110101010001010110010",
"110110101000101101011101",
"110110100111010000001110",
"110110100101110011000011",
"110110100100010101111101",
"110110100010111000111100",
"110110100001011100000000",
"110110011111111111001010",
"110110011110100010011000",
"110110011101000101101010",
"110110011011101001000010",
"110110011010001100011111",
"110110011000110000000001",
"110110010111010011100111",
"110110010101110111010011",
"110110010100011011000011",
"110110010010111110111001",
"110110010001100010110011",
"110110010000000110110010",
"110110001110101010110110",
"110110001101001110111111",
"110110001011110011001100",
"110110001010010111011111",
"110110001000111011110110",
"110110000111100000010011",
"110110000110000100110100",
"110110000100101001011010",
"110110000011001110000100",
"110110000001110010110100",
"110110000000010111101000",
"110101111110111100100001",
"110101111101100001011111",
"110101111100000110100010",
"110101111010101011101010",
"110101111001010000110110",
"110101110111110110000111",
"110101110110011011011101",
"110101110101000000111000",
"110101110011100110010111",
"110101110010001011111011",
"110101110000110001100100",
"110101101111010111010010",
"110101101101111101000100",
"110101101100100010111011",
"110101101011001000110111",
"110101101001101110110111",
"110101101000010100111101",
"110101100110111011000111",
"110101100101100001010101",
"110101100100000111101001",
"110101100010101110000001",
"110101100001010100011110",
"110101011111111010111111",
"110101011110100001100101",
"110101011101001000010000",
"110101011011101110111111",
"110101011010010101110011",
"110101011000111100101100",
"110101010111100011101001",
"110101010110001010101100",
"110101010100110001110010",
"110101010011011000111101",
"110101010010000000001101",
"110101010000100111100010",
"110101001111001110111011",
"110101001101110110011001",
"110101001100011101111011",
"110101001011000101100010",
"110101001001101101001101",
"110101001000010100111110",
"110101000110111100110010",
"110101000101100100101011",
"110101000100001100101001",
"110101000010110100101100",
"110101000001011100110011",
"110101000000000100111110",
"110100111110101101001110",
"110100111101010101100011",
"110100111011111101111100",
"110100111010100110011001",
"110100111001001110111011",
"110100110111110111100010",
"110100110110100000001101",
"110100110101001000111101",
"110100110011110001110001",
"110100110010011010101010",
"110100110001000011100111",
"110100101111101100101000",
"110100101110010101101111",
"110100101100111110111001",
"110100101011101000001000",
"110100101010010001011100",
"110100101000111010110100",
"110100100111100100010000",
"110100100110001101110001",
"110100100100110111010110",
"110100100011100001000000",
"110100100010001010101110",
"110100100000110100100001",
"110100011111011110011000",
"110100011110001000010011",
"110100011100110010010011",
"110100011011011100010111",
"110100011010000110100000",
"110100011000110000101101",
"110100010111011010111110",
"110100010110000101010100",
"110100010100101111101110",
"110100010011011010001101",
"110100010010000100110000",
"110100010000101111010111",
"110100001111011010000011",
"110100001110000100110011",
"110100001100101111100111",
"110100001011011010100000",
"110100001010000101011101",
"110100001000110000011110",
"110100000111011011100100",
"110100000110000110101110",
"110100000100110001111100",
"110100000011011101001111",
"110100000010001000100110",
"110100000000110100000001",
"110011111111011111100000",
"110011111110001011000100",
"110011111100110110101100",
"110011111011100010011001",
"110011111010001110001001",
"110011111000111001111110",
"110011110111100101110111",
"110011110110010001110101",
"110011110100111101110110",
"110011110011101001111100",
"110011110010010110000110",
"110011110001000010010101",
"110011101111101110100111",
"110011101110011010111110",
"110011101101000111011001",
"110011101011110011111001",
"110011101010100000011100",
"110011101001001101000100",
"110011100111111001110000",
"110011100110100110100000",
"110011100101010011010100",
"110011100100000000001101",
"110011100010101101001010",
"110011100001011010001010",
"110011100000000111010000",
"110011011110110100011001",
"110011011101100001100110",
"110011011100001110111000",
"110011011010111100001101",
"110011011001101001100111",
"110011011000010111000101",
"110011010111000100100111",
"110011010101110010001110",
"110011010100011111111000",
"110011010011001101100111",
"110011010001111011011001",
"110011010000101001010000",
"110011001111010111001011",
"110011001110000101001010",
"110011001100110011001101",
"110011001011100001010100",
"110011001010001111011111",
"110011001000111101101111",
"110011000111101100000010",
"110011000110011010011010",
"110011000101001000110101",
"110011000011110111010101",
"110011000010100101111000",
"110011000001010100100000",
"110011000000000011001100",
"110010111110110001111100",
"110010111101100000110000",
"110010111100001111101000",
"110010111010111110100100",
"110010111001101101100100",
"110010111000011100101000",
"110010110111001011110000",
"110010110101111010111100",
"110010110100101010001100",
"110010110011011001100000",
"110010110010001000111000",
"110010110000111000010100",
"110010101111100111110100",
"110010101110010111011000",
"110010101101000111000000",
"110010101011110110101100",
"110010101010100110011100",
"110010101001010110010000",
"110010101000000110001000",
"110010100110110110000100",
"110010100101100110000100",
"110010100100010110001000",
"110010100011000110010000",
"110010100001110110011011",
"110010100000100110101011",
"110010011111010110111111",
"110010011110000111010110",
"110010011100110111110001",
"110010011011101000010001",
"110010011010011000110100",
"110010011001001001011011",
"110010010111111010000110",
"110010010110101010110101",
"110010010101011011101000",
"110010010100001100011111",
"110010010010111101011001",
"110010010001101110011000",
"110010010000011111011010",
"110010001111010000100001",
"110010001110000001101011",
"110010001100110010111001",
"110010001011100100001011",
"110010001010010101100000",
"110010001001000110111010",
"110010000111111000010111",
"110010000110101001111001",
"110010000101011011011110",
"110010000100001101000111",
"110010000010111110110011",
"110010000001110000100100",
"110010000000100010011000",
"110001111111010100010001",
"110001111110000110001101",
"110001111100111000001100",
"110001111011101010010000",
"110001111010011100011000",
"110001111001001110100011",
"110001111000000000110010",
"110001110110110011000101",
"110001110101100101011011",
"110001110100010111110110",
"110001110011001010010100",
"110001110001111100110110",
"110001110000101111011011",
"110001101111100010000101",
"110001101110010100110010",
"110001101101000111100011",
"110001101011111010011000",
"110001101010101101010000",
"110001101001100000001100",
"110001101000010011001100",
"110001100111000110010000",
"110001100101111001010111",
"110001100100101100100010",
"110001100011011111110001",
"110001100010010011000100",
"110001100001000110011010",
"110001011111111001110100",
"110001011110101101010010",
"110001011101100000110011",
"110001011100010100011000",
"110001011011001000000001",
"110001011001111011101101",
"110001011000101111011101",
"110001010111100011010001",
"110001010110010111001000",
"110001010101001011000100",
"110001010011111111000010",
"110001010010110011000101",
"110001010001100111001011",
"110001010000011011010101",
"110001001111001111100010",
"110001001110000011110011",
"110001001100111000001000",
"110001001011101100100000",
"110001001010100000111100",
"110001001001010101011011",
"110001001000001001111111",
"110001000110111110100101",
"110001000101110011010000",
"110001000100100111111110",
"110001000011011100110000",
"110001000010010001100101",
"110001000001000110011110",
"110000111111111011011010",
"110000111110110000011010",
"110000111101100101011110",
"110000111100011010100101",
"110000111011001111110000",
"110000111010000100111110",
"110000111000111010010000",
"110000110111101111100101",
"110000110110100100111110",
"110000110101011010011011",
"110000110100001111111011",
"110000110011000101011111",
"110000110001111011000110",
"110000110000110000110001",
"110000101111100110011111",
"110000101110011100010001",
"110000101101010010000110",
"110000101100000111111111",
"110000101010111101111100",
"110000101001110011111100",
"110000101000101001111111",
"110000100111100000000110",
"110000100110010110010001",
"110000100101001100011111",
"110000100100000010110000",
"110000100010111001000101",
"110000100001101111011110",
"110000100000100101111001",
"110000011111011100011001",
"110000011110010010111100",
"110000011101001001100010",
"110000011100000000001100",
"110000011010110110111001",
"110000011001101101101010",
"110000011000100100011111",
"110000010111011011010110",
"110000010110010010010001",
"110000010101001001010000",
"110000010100000000010010",
"110000010010110111011000",
"110000010001101110100001",
"110000010000100101101101",
"110000001111011100111101",
"110000001110010100010000",
"110000001101001011100111",
"110000001100000011000001",
"110000001010111010011110",
"110000001001110001111111",
"110000001000101001100011",
"110000000111100001001011",
"110000000110011000110110",
"110000000101010000100101",
"110000000100001000010111",
"110000000011000000001100",
"110000000001111000000101",
"110000000000110000000001",
"101111111111101000000000",
"101111111110100000000011",
"101111111101011000001001",
"101111111100010000010011",
"101111111011001000100000",
"101111111010000000110000",
"101111111000111001000100",
"101111110111110001011011",
"101111110110101001110101",
"101111110101100010010010",
"101111110100011010110100",
"101111110011010011011000",
"101111110010001100000000",
"101111110001000100101011",
"101111101111111101011001",
"101111101110110110001011",
"101111101101101111000000",
"101111101100100111111000",
"101111101011100000110011",
"101111101010011001110010",
"101111101001010010110101",
"101111101000001011111010",
"101111100111000101000011",
"101111100101111110001111",
"101111100100110111011110",
"101111100011110000110001",
"101111100010101010000111",
"101111100001100011100000",
"101111100000011100111101",
"101111011111010110011101",
"101111011110010000000000",
"101111011101001001100110",
"101111011100000011010000",
"101111011010111100111100",
"101111011001110110101100",
"101111011000110000100000",
"101111010111101010010110",
"101111010110100100010000",
"101111010101011110001101",
"101111010100011000001110",
"101111010011010010010001",
"101111010010001100011000",
"101111010001000110100010",
"101111010000000000101111",
"101111001110111011000000",
"101111001101110101010011",
"101111001100101111101010",
"101111001011101010000100",
"101111001010100100100010",
"101111001001011111000010",
"101111001000011001100110",
"101111000111010100001101",
"101111000110001110110111",
"101111000101001001100100",
"101111000100000100010100",
"101111000010111111001000",
"101111000001111001111111",
"101111000000110100111001",
"101110111111101111110110",
"101110111110101010110110",
"101110111101100101111010",
"101110111100100001000001",
"101110111011011100001010",
"101110111010010111010111",
"101110111001010010100111",
"101110111000001101111011",
"101110110111001001010001",
"101110110110000100101011",
"101110110101000000000111",
"101110110011111011100111",
"101110110010110111001010",
"101110110001110010110000",
"101110110000101110011001",
"101110101111101010000110",
"101110101110100101110101",
"101110101101100001101000",
"101110101100011101011101",
"101110101011011001010110",
"101110101010010101010010",
"101110101001010001010001",
"101110101000001101010011",
"101110100111001001011000",
"101110100110000101100000",
"101110100101000001101100",
"101110100011111101111010",
"101110100010111010001100",
"101110100001110110100000",
"101110100000110010111000",
"101110011111101111010011",
"101110011110101011110000",
"101110011101101000010001",
"101110011100100100110101",
"101110011011100001011100",
"101110011010011110000110",
"101110011001011010110011",
"101110011000010111100011",
"101110010111010100010111",
"101110010110010001001101",
"101110010101001110000110",
"101110010100001011000010",
"101110010011001000000010",
"101110010010000101000100",
"101110010001000010001001",
"101110001111111111010010",
"101110001110111100011101",
"101110001101111001101100",
"101110001100110110111101",
"101110001011110100010001",
"101110001010110001101001",
"101110001001101111000011",
"101110001000101100100001",
"101110000111101010000001",
"101110000110100111100101",
"101110000101100101001011",
"101110000100100010110101",
"101110000011100000100001",
"101110000010011110010001",
"101110000001011100000011",
"101110000000011001111000",
"101101111111010111110001",
"101101111110010101101100",
"101101111101010011101010",
"101101111100010001101011",
"101101111011001111101111",
"101101111010001101110111",
"101101111001001100000001",
"101101111000001010001110",
"101101110111001000011110",
"101101110110000110110001",
"101101110101000101000111",
"101101110100000011011111",
"101101110011000001111011",
"101101110010000000011010",
"101101110000111110111011",
"101101101111111101100000",
"101101101110111100000111",
"101101101101111010110010",
"101101101100111001011111",
"101101101011111000001111",
"101101101010110111000010",
"101101101001110101111000",
"101101101000110100110001",
"101101100111110011101101",
"101101100110110010101100",
"101101100101110001101101",
"101101100100110000110010",
"101101100011101111111001",
"101101100010101111000100",
"101101100001101110010001",
"101101100000101101100001",
"101101011111101100110100",
"101101011110101100001001",
"101101011101101011100010",
"101101011100101010111110",
"101101011011101010011100",
"101101011010101001111101",
"101101011001101001100001",
"101101011000101001001000",
"101101010111101000110010",
"101101010110101000011111",
"101101010101101000001110",
"101101010100101000000001",
"101101010011100111110110",
"101101010010100111101110",
"101101010001100111101001",
"101101010000100111100111",
"101101001111100111100111",
"101101001110100111101010",
"101101001101100111110001",
"101101001100100111111010",
"101101001011101000000101",
"101101001010101000010100",
"101101001001101000100110",
"101101001000101000111010",
"101101000111101001010001",
"101101000110101001101011",
"101101000101101010000111",
"101101000100101010100111",
"101101000011101011001001",
"101101000010101011101110",
"101101000001101100010110",
"101101000000101101000001",
"101100111111101101101110",
"101100111110101110011110",
"101100111101101111010001",
"101100111100110000000111",
"101100111011110001000000",
"101100111010110001111011",
"101100111001110010111001",
"101100111000110011111010",
"101100110111110100111101",
"101100110110110110000100",
"101100110101110111001101",
"101100110100111000011001",
"101100110011111001100111",
"101100110010111010111000",
"101100110001111100001101",
"101100110000111101100011",
"101100101111111110111101",
"101100101111000000011001",
"101100101110000001111000",
"101100101101000011011010",
"101100101100000100111110",
"101100101011000110100110",
"101100101010001000010000",
"101100101001001001111100",
"101100101000001011101100",
"101100100111001101011110",
"101100100110001111010010",
"101100100101010001001010",
"101100100100010011000100",
"101100100011010101000001",
"101100100010010111000001",
"101100100001011001000011",
"101100100000011011001000",
"101100011111011101001111",
"101100011110011111011010",
"101100011101100001100111",
"101100011100100011110111",
"101100011011100110001001",
"101100011010101000011110",
"101100011001101010110110",
"101100011000101101010000",
"101100010111101111101101",
"101100010110110010001101",
"101100010101110100101111",
"101100010100110111010101",
"101100010011111001111100",
"101100010010111100100111",
"101100010001111111010100",
"101100010001000010000011",
"101100010000000100110110",
"101100001111000111101011",
"101100001110001010100010",
"101100001101001101011101",
"101100001100010000011010",
"101100001011010011011001",
"101100001010010110011011",
"101100001001011001100000",
"101100001000011100100111",
"101100000111011111110010",
"101100000110100010111110",
"101100000101100110001101",
"101100000100101001011111",
"101100000011101100110100",
"101100000010110000001011",
"101100000001110011100101",
"101100000000110111000001",
"101011111111111010100000",
"101011111110111110000010",
"101011111110000001100110",
"101011111101000101001100",
"101011111100001000110110",
"101011111011001100100010",
"101011111010010000010000",
"101011111001010100000001",
"101011111000010111110101",
"101011110111011011101011",
"101011110110011111100100",
"101011110101100011011111",
"101011110100100111011101",
"101011110011101011011110",
"101011110010101111100001",
"101011110001110011100111",
"101011110000110111101111",
"101011101111111011111010",
"101011101111000000000111",
"101011101110000100010111",
"101011101101001000101001",
"101011101100001100111110",
"101011101011010001010110",
"101011101010010101110000",
"101011101001011010001100",
"101011101000011110101011",
"101011100111100011001101",
"101011100110100111110001",
"101011100101101100011000",
"101011100100110001000001",
"101011100011110101101101",
"101011100010111010011011",
"101011100001111111001100",
"101011100001000100000000",
"101011100000001000110110",
"101011011111001101101110",
"101011011110010010101001",
"101011011101010111100110",
"101011011100011100100110",
"101011011011100001101001",
"101011011010100110101101",
"101011011001101011110101",
"101011011000110000111111",
"101011010111110110001011",
"101011010110111011011010",
"101011010110000000101011",
"101011010101000101111111",
"101011010100001011010110",
"101011010011010000101110",
"101011010010010110001010",
"101011010001011011100111",
"101011010000100001001000",
"101011001111100110101010",
"101011001110101100010000",
"101011001101110001110111",
"101011001100110111100001",
"101011001011111101001110",
"101011001011000010111101",
"101011001010001000101110",
"101011001001001110100010",
"101011001000010100011001",
"101011000111011010010010",
"101011000110100000001101",
"101011000101100110001011",
"101011000100101100001011",
"101011000011110010001101",
"101011000010111000010010",
"101011000001111110011010",
"101011000001000100100100",
"101011000000001010110000",
"101010111111010000111111",
"101010111110010111010000",
"101010111101011101100100",
"101010111100100011111010",
"101010111011101010010010",
"101010111010110000101101",
"101010111001110111001010",
"101010111000111101101010",
"101010111000000100001100",
"101010110111001010110000",
"101010110110010001010111",
"101010110101011000000001",
"101010110100011110101100",
"101010110011100101011010",
"101010110010101100001011",
"101010110001110010111110",
"101010110000111001110011",
"101010110000000000101011",
"101010101111000111100101",
"101010101110001110100001",
"101010101101010101100000",
"101010101100011100100001",
"101010101011100011100101",
"101010101010101010101011",
"101010101001110001110011",
"101010101000111000111110",
"101010101000000000001011",
"101010100111000111011010",
"101010100110001110101100",
"101010100101010110000000",
"101010100100011101010110",
"101010100011100100101111",
"101010100010101100001010",
"101010100001110011101000",
"101010100000111011001000",
"101010100000000010101010",
"101010011111001010001111",
"101010011110010001110101",
"101010011101011001011111",
"101010011100100001001010",
"101010011011101000111000",
"101010011010110000101000",
"101010011001111000011011",
"101010011001000000010000",
"101010011000001000000111",
"101010010111010000000001",
"101010010110010111111101",
"101010010101011111111011",
"101010010100100111111011",
"101010010011101111111110",
"101010010010111000000011",
"101010010010000000001011",
"101010010001001000010100",
"101010010000010000100000",
"101010001111011000101111",
"101010001110100000111111",
"101010001101101001010010",
"101010001100110001101000",
"101010001011111001111111",
"101010001011000010011001",
"101010001010001010110101",
"101010001001010011010011",
"101010001000011011110100",
"101010000111100100010111",
"101010000110101100111100",
"101010000101110101100100",
"101010000100111110001110",
"101010000100000110111010",
"101010000011001111101000",
"101010000010011000011001",
"101010000001100001001100",
"101010000000101010000001",
"101001111111110010111000",
"101001111110111011110010",
"101001111110000100101110",
"101001111101001101101100",
"101001111100010110101100",
"101001111011011111101111",
"101001111010101000110100",
"101001111001110001111011",
"101001111000111011000101",
"101001111000000100010000",
"101001110111001101011110",
"101001110110010110101110",
"101001110101100000000001",
"101001110100101001010101",
"101001110011110010101100",
"101001110010111100000101",
"101001110010000101100001",
"101001110001001110111110",
"101001110000011000011110",
"101001101111100010000000",
"101001101110101011100100",
"101001101101110101001010",
"101001101100111110110011",
"101001101100001000011110",
"101001101011010010001011",
"101001101010011011111010",
"101001101001100101101100",
"101001101000101111011111",
"101001100111111001010101",
"101001100111000011001101",
"101001100110001101001000",
"101001100101010111000100",
"101001100100100001000011",
"101001100011101011000100",
"101001100010110101000111",
"101001100001111111001100",
"101001100001001001010100",
"101001100000010011011101",
"101001011111011101101001",
"101001011110100111110111",
"101001011101110010000111",
"101001011100111100011001",
"101001011100000110101110",
"101001011011010001000101",
"101001011010011011011101",
"101001011001100101111000",
"101001011000110000010110",
"101001010111111010110101",
"101001010111000101010111",
"101001010110001111111010",
"101001010101011010100000",
"101001010100100101001000",
"101001010011101111110010",
"101001010010111010011110",
"101001010010000101001101",
"101001010001001111111101",
"101001010000011010110000",
"101001001111100101100101",
"101001001110110000011100",
"101001001101111011010101",
"101001001101000110010000",
"101001001100010001001110",
"101001001011011100001101",
"101001001010100111001111",
"101001001001110010010011",
"101001001000111101011001",
"101001001000001000100001",
"101001000111010011101011",
"101001000110011110110111",
"101001000101101010000110",
"101001000100110101010110",
"101001000100000000101001",
"101001000011001011111110",
"101001000010010111010101",
"101001000001100010101110",
"101001000000101110001001",
"101000111111111001100110",
"101000111111000101000101",
"101000111110010000100111",
"101000111101011100001010",
"101000111100100111110000",
"101000111011110011011000",
"101000111010111111000001",
"101000111010001010101101",
"101000111001010110011011",
"101000111000100010001011",
"101000110111101101111101",
"101000110110111001110010",
"101000110110000101101000",
"101000110101010001100000",
"101000110100011101011011",
"101000110011101001010111",
"101000110010110101010110",
"101000110010000001010111",
"101000110001001101011001",
"101000110000011001011110",
"101000101111100101100101",
"101000101110110001101110",
"101000101101111101111001",
"101000101101001010000110",
"101000101100010110010101",
"101000101011100010100111",
"101000101010101110111010",
"101000101001111011001111",
"101000101001000111100110",
"101000101000010100000000",
"101000100111100000011011",
"101000100110101100111001",
"101000100101111001011000",
"101000100101000101111010",
"101000100100010010011110",
"101000100011011111000011",
"101000100010101011101011",
"101000100001111000010101",
"101000100001000101000000",
"101000100000010001101110",
"101000011111011110011110",
"101000011110101011010000",
"101000011101111000000100",
"101000011101000100111010",
"101000011100010001110001",
"101000011011011110101011",
"101000011010101011100111",
"101000011001111000100101",
"101000011001000101100101",
"101000011000010010100111",
"101000010111011111101011",
"101000010110101100110001",
"101000010101111001111001",
"101000010101000111000011",
"101000010100010100001111",
"101000010011100001011101",
"101000010010101110101101",
"101000010001111011111111",
"101000010001001001010011",
"101000010000010110101001",
"101000001111100100000001",
"101000001110110001011011",
"101000001101111110110111",
"101000001101001100010101",
"101000001100011001110101",
"101000001011100111010111",
"101000001010110100111011",
"101000001010000010100001",
"101000001001010000001000",
"101000001000011101110010",
"101000000111101011011110",
"101000000110111001001100",
"101000000110000110111100",
"101000000101010100101101",
"101000000100100010100001",
"101000000011110000010111",
"101000000010111110001110",
"101000000010001100001000",
"101000000001011010000011",
"101000000000101000000001",
"100111111111110110000000",
"100111111111000100000001",
"100111111110010010000101",
"100111111101100000001010",
"100111111100101110010001",
"100111111011111100011010",
"100111111011001010100101",
"100111111010011000110011",
"100111111001100111000010",
"100111111000110101010010",
"100111111000000011100101",
"100111110111010001111010",
"100111110110100000010001",
"100111110101101110101001",
"100111110100111101000100",
"100111110100001011100001",
"100111110011011001111111",
"100111110010101000011111",
"100111110001110111000010",
"100111110001000101100110",
"100111110000010100001100",
"100111101111100010110100",
"100111101110110001011110",
"100111101110000000001010",
"100111101101001110111000",
"100111101100011101100111",
"100111101011101100011001",
"100111101010111011001101",
"100111101010001010000010",
"100111101001011000111001",
"100111101000100111110011",
"100111100111110110101110",
"100111100111000101101011",
"100111100110010100101010",
"100111100101100011101010",
"100111100100110010101101",
"100111100100000001110010",
"100111100011010000111000",
"100111100010100000000001",
"100111100001101111001011",
"100111100000111110010111",
"100111100000001101100101",
"100111011111011100110101",
"100111011110101100000111",
"100111011101111011011010",
"100111011101001010110000",
"100111011100011010000111",
"100111011011101001100001",
"100111011010111000111100",
"100111011010001000011001",
"100111011001010111111000",
"100111011000100111011001",
"100111010111110110111011",
"100111010111000110100000",
"100111010110010110000110",
"100111010101100101101110",
"100111010100110101011000",
"100111010100000101000100",
"100111010011010100110010",
"100111010010100100100010",
"100111010001110100010011",
"100111010001000100000111",
"100111010000010011111100",
"100111001111100011110011",
"100111001110110011101100",
"100111001110000011100110",
"100111001101010011100011",
"100111001100100011100001",
"100111001011110011100010",
"100111001011000011100100",
"100111001010010011101000",
"100111001001100011101101",
"100111001000110011110101",
"100111001000000011111110",
"100111000111010100001010",
"100111000110100100010111",
"100111000101110100100101",
"100111000101000100110110",
"100111000100010101001001",
"100111000011100101011101",
"100111000010110101110011",
"100111000010000110001011",
"100111000001010110100101",
"100111000000100111000001",
"100110111111110111011110",
"100110111111000111111101",
"100110111110011000011110",
"100110111101101001000001",
"100110111100111001100110",
"100110111100001010001100",
"100110111011011010110101",
"100110111010101011011111",
"100110111001111100001010",
"100110111001001100111000",
"100110111000011101101000",
"100110110111101110011001",
"100110110110111111001100",
"100110110110010000000001",
"100110110101100000110111",
"100110110100110001110000",
"100110110100000010101010",
"100110110011010011100110",
"100110110010100100100100",
"100110110001110101100011",
"100110110001000110100100",
"100110110000010111100111",
"100110101111101000101100",
"100110101110111001110011",
"100110101110001010111011",
"100110101101011100000110",
"100110101100101101010010",
"100110101011111110011111",
"100110101011001111101111",
"100110101010100001000000",
"100110101001110010010011",
"100110101001000011101000",
"100110101000010100111110",
"100110100111100110010111",
"100110100110110111110001",
"100110100110001001001101",
"100110100101011010101010",
"100110100100101100001001",
"100110100011111101101011",
"100110100011001111001101",
"100110100010100000110010",
"100110100001110010011000",
"100110100001000100000000",
"100110100000010101101010",
"100110011111100111010110",
"100110011110111001000011",
"100110011110001010110010",
"100110011101011100100011",
"100110011100101110010101",
"100110011100000000001010",
"100110011011010010000000",
"100110011010100011110111",
"100110011001110101110001",
"100110011001000111101100",
"100110011000011001101001",
"100110010111101011100111",
"100110010110111101101000",
"100110010110001111101010",
"100110010101100001101110",
"100110010100110011110011",
"100110010100000101111010",
"100110010011011000000011",
"100110010010101010001110",
"100110010001111100011010",
"100110010001001110101000",
"100110010000100000111000",
"100110001111110011001010",
"100110001111000101011101",
"100110001110010111110010",
"100110001101101010001000",
"100110001100111100100001",
"100110001100001110111011",
"100110001011100001010111",
"100110001010110011110100",
"100110001010000110010011",
"100110001001011000110100",
"100110001000101011010110",
"100110000111111101111011",
"100110000111010000100000",
"100110000110100011001000",
"100110000101110101110001",
"100110000101001000011100",
"100110000100011011001001",
"100110000011101101110111",
"100110000011000000100111",
"100110000010010011011001",
"100110000001100110001100",
"100110000000111001000001",
"100110000000001011111000",
"100101111111011110110000",
"100101111110110001101011",
"100101111110000100100110",
"100101111101010111100100",
"100101111100101010100011",
"100101111011111101100100",
"100101111011010000100110",
"100101111010100011101010",
"100101111001110110110000",
"100101111001001001110111",
"100101111000011101000000",
"100101110111110000001011",
"100101110111000011010111",
"100101110110010110100101",
"100101110101101001110101",
"100101110100111101000110",
"100101110100010000011001",
"100101110011100011101110",
"100101110010110111000100",
"100101110010001010011100",
"100101110001011101110110",
"100101110000110001010001",
"100101110000000100101110",
"100101101111011000001101",
"100101101110101011101101",
"100101101101111111001110",
"100101101101010010110010",
"100101101100100110010111",
"100101101011111001111110",
"100101101011001101100110",
"100101101010100001010000",
"100101101001110100111100",
"100101101001001000101001",
"100101101000011100011000",
"100101100111110000001000",
"100101100111000011111010",
"100101100110010111101110",
"100101100101101011100011",
"100101100100111111011010",
"100101100100010011010011",
"100101100011100111001101",
"100101100010111011001001",
"100101100010001111000111",
"100101100001100011000110",
"100101100000110111000110",
"100101100000001011001001",
"100101011111011111001100",
"100101011110110011010010",
"100101011110000111011001",
"100101011101011011100010",
"100101011100101111101100",
"100101011100000011111000",
"100101011011011000000110",
"100101011010101100010101",
"100101011010000000100101",
"100101011001010100111000",
"100101011000101001001100",
"100101010111111101100001",
"100101010111010001111000",
"100101010110100110010001",
"100101010101111010101011",
"100101010101001111000111",
"100101010100100011100101",
"100101010011111000000100",
"100101010011001100100100",
"100101010010100001000111",
"100101010001110101101010",
"100101010001001010010000",
"100101010000011110110111",
"100101001111110011011111",
"100101001111001000001001",
"100101001110011100110101",
"100101001101110001100010",
"100101001101000110010001",
"100101001100011011000010",
"100101001011101111110100",
"100101001011000100100111",
"100101001010011001011100",
"100101001001101110010011",
"100101001001000011001011",
"100101001000011000000101",
"100101000111101101000000",
"100101000111000001111101",
"100101000110010110111100",
"100101000101101011111100",
"100101000101000000111101",
"100101000100010110000001",
"100101000011101011000101",
"100101000011000000001100",
"100101000010010101010011",
"100101000001101010011101",
"100101000000111111101000",
"100101000000010100110100",
"100100111111101010000010",
"100100111110111111010010",
"100100111110010100100011",
"100100111101101001110110",
"100100111100111111001010",
"100100111100010100011111",
"100100111011101001110111",
"100100111010111111010000",
"100100111010010100101010",
"100100111001101010000110",
"100100111000111111100011",
"100100111000010101000010",
"100100110111101010100011",
"100100110111000000000101",
"100100110110010101101000",
"100100110101101011001101",
"100100110101000000110100",
"100100110100010110011100",
"100100110011101100000110",
"100100110011000001110001",
"100100110010010111011101",
"100100110001101101001100",
"100100110001000010111011",
"100100110000011000101101",
"100100101111101110011111",
"100100101111000100010100",
"100100101110011010001001",
"100100101101110000000001",
"100100101101000101111001",
"100100101100011011110100",
"100100101011110001101111",
"100100101011000111101101",
"100100101010011101101100",
"100100101001110011101100",
"100100101001001001101110",
"100100101000011111110001",
"100100100111110101110110",
"100100100111001011111100",
"100100100110100010000100",
"100100100101111000001101",
"100100100101001110011000",
"100100100100100100100101",
"100100100011111010110010",
"100100100011010001000010",
"100100100010100111010010",
"100100100001111101100101",
"100100100001010011111001",
"100100100000101010001110",
"100100100000000000100101",
"100100011111010110111101",
"100100011110101101010110",
"100100011110000011110010",
"100100011101011010001110",
"100100011100110000101100",
"100100011100000111001100",
"100100011011011101101101",
"100100011010110100010000",
"100100011010001010110100",
"100100011001100001011001",
"100100011000111000000000",
"100100011000001110101001",
"100100010111100101010011",
"100100010110111011111110",
"100100010110010010101011",
"100100010101101001011001",
"100100010101000000001001",
"100100010100010110111010",
"100100010011101101101101",
"100100010011000100100001",
"100100010010011011010111",
"100100010001110010001110",
"100100010001001001000111",
"100100010000100000000001",
"100100001111110110111100",
"100100001111001101111001",
"100100001110100100110111",
"100100001101111011110111",
"100100001101010010111000",
"100100001100101001111011",
"100100001100000000111111",
"100100001011011000000101",
"100100001010101111001100",
"100100001010000110010101",
"100100001001011101011110",
"100100001000110100101010",
"100100001000001011110111",
"100100000111100011000101",
"100100000110111010010101",
"100100000110010001100110",
"100100000101101000111000",
"100100000101000000001100",
"100100000100010111100010",
"100100000011101110111001",
"100100000011000110010001",
"100100000010011101101011",
"100100000001110101000110",
"100100000001001100100011",
"100100000000100100000001",
"100011111111111011100000",
"100011111111010011000001",
"100011111110101010100011",
"100011111110000010000111",
"100011111101011001101100",
"100011111100110001010011",
"100011111100001000111011",
"100011111011100000100100",
"100011111010111000001111",
"100011111010001111111011",
"100011111001100111101001",
"100011111000111111011000",
"100011111000010111001000",
"100011110111101110111010",
"100011110111000110101101",
"100011110110011110100010",
"100011110101110110011000",
"100011110101001110001111",
"100011110100100110001000",
"100011110011111110000011",
"100011110011010101111110",
"100011110010101101111011",
"100011110010000101111010",
"100011110001011101111010",
"100011110000110101111011",
"100011110000001101111110",
"100011101111100110000010",
"100011101110111110000111",
"100011101110010110001110",
"100011101101101110010111",
"100011101101000110100000",
"100011101100011110101011",
"100011101011110110111000",
"100011101011001111000101",
"100011101010100111010101",
"100011101001111111100101",
"100011101001010111110111",
"100011101000110000001011",
"100011101000001000011111",
"100011100111100000110101",
"100011100110111001001101",
"100011100110010001100110",
"100011100101101010000000",
"100011100101000010011100",
"100011100100011010111001",
"100011100011110011010111",
"100011100011001011110111",
"100011100010100100011000",
"100011100001111100111010",
"100011100001010101011110",
"100011100000101110000011",
"100011100000000110101010",
"100011011111011111010010",
"100011011110110111111011",
"100011011110010000100110",
"100011011101101001010010",
"100011011101000001111111",
"100011011100011010101110",
"100011011011110011011110",
"100011011011001100010000",
"100011011010100101000011",
"100011011001111101110111",
"100011011001010110101100",
"100011011000101111100011",
"100011011000001000011100",
"100011010111100001010101",
"100011010110111010010000",
"100011010110010011001100",
"100011010101101100001010",
"100011010101000101001001",
"100011010100011110001001",
"100011010011110111001011",
"100011010011010000001110",
"100011010010101001010010",
"100011010010000010011000",
"100011010001011011011111",
"100011010000110100101000",
"100011010000001101110001",
"100011001111100110111100",
"100011001111000000001001",
"100011001110011001010111",
"100011001101110010100110",
"100011001101001011110110",
"100011001100100101001000",
"100011001011111110011011",
"100011001011010111101111",
"100011001010110001000101",
"100011001010001010011100",
"100011001001100011110100",
"100011001000111101001110",
"100011001000010110101001",
"100011000111110000000101",
"100011000111001001100011",
"100011000110100011000010",
"100011000101111100100010",
"100011000101010110000100",
"100011000100101111100111",
"100011000100001001001011",
"100011000011100010110001",
"100011000010111100011000",
"100011000010010110000000",
"100011000001101111101010",
"100011000001001001010100",
"100011000000100011000001",
"100010111111111100101110",
"100010111111010110011101",
"100010111110110000001101",
"100010111110001001111110",
"100010111101100011110001",
"100010111100111101100101",
"100010111100010111011010",
"100010111011110001010001",
"100010111011001011001001",
"100010111010100101000010",
"100010111001111110111100",
"100010111001011000111000",
"100010111000110010110101",
"100010111000001100110100",
"100010110111100110110011",
"100010110111000000110100",
"100010110110011010110111",
"100010110101110100111010",
"100010110101001110111111",
"100010110100101001000101",
"100010110100000011001101",
"100010110011011101010101",
"100010110010110111011111",
"100010110010010001101011",
"100010110001101011110111",
"100010110001000110000101",
"100010110000100000010100",
"100010101111111010100101",
"100010101111010100110110",
"100010101110101111001001",
"100010101110001001011101",
"100010101101100011110011",
"100010101100111110001010",
"100010101100011000100010",
"100010101011110010111011",
"100010101011001101010110",
"100010101010100111110010",
"100010101010000010001111",
"100010101001011100101101",
"100010101000110111001101",
"100010101000010001101110",
"100010100111101100010000",
"100010100111000110110100",
"100010100110100001011001",
"100010100101111011111111",
"100010100101010110100110",
"100010100100110001001111",
"100010100100001011111000",
"100010100011100110100100",
"100010100011000001010000",
"100010100010011011111110",
"100010100001110110101100",
"100010100001010001011101",
"100010100000101100001110",
"100010100000000111000001",
"100010011111100001110100",
"100010011110111100101010",
"100010011110010111100000",
"100010011101110010011000",
"100010011101001101010000",
"100010011100101000001011",
"100010011100000011000110",
"100010011011011110000011",
"100010011010111001000001",
"100010011010010100000000",
"100010011001101111000000",
"100010011001001010000010",
"100010011000100101000100",
"100010011000000000001001",
"100010010111011011001110",
"100010010110110110010101",
"100010010110010001011100",
"100010010101101100100101",
"100010010101000111110000",
"100010010100100010111011",
"100010010011111110001000",
"100010010011011001010110",
"100010010010110100100101",
"100010010010001111110110",
"100010010001101011000111",
"100010010001000110011010",
"100010010000100001101110",
"100010001111111101000100",
"100010001111011000011010",
"100010001110110011110010",
"100010001110001111001011",
"100010001101101010100101",
"100010001101000110000001",
"100010001100100001011110",
"100010001011111100111011",
"100010001011011000011011",
"100010001010110011111011",
"100010001010001111011101",
"100010001001101010111111",
"100010001001000110100011",
"100010001000100010001001",
"100010000111111101101111",
"100010000111011001010111",
"100010000110110100111111",
"100010000110010000101010",
"100010000101101100010101",
"100010000101001000000001",
"100010000100100011101111",
"100010000011111111011110",
"100010000011011011001110",
"100010000010110110111111",
"100010000010010010110010",
"100010000001101110100110",
"100010000001001010011011",
"100010000000100110010001",
"100010000000000010001000",
"100001111111011110000001",
"100001111110111001111010",
"100001111110010101110101",
"100001111101110001110001",
"100001111101001101101111",
"100001111100101001101101",
"100001111100000101101101",
"100001111011100001101110",
"100001111010111101110000",
"100001111010011001110011",
"100001111001110101111000",
"100001111001010001111101",
"100001111000101110000100",
"100001111000001010001100",
"100001110111100110010101",
"100001110111000010100000",
"100001110110011110101011",
"100001110101111010111000",
"100001110101010111000110",
"100001110100110011010101",
"100001110100001111100110",
"100001110011101011110111",
"100001110011001000001010",
"100001110010100100011110",
"100001110010000000110011",
"100001110001011101001001",
"100001110000111001100000",
"100001110000010101111001",
"100001101111110010010011",
"100001101111001110101110",
"100001101110101011001010",
"100001101110000111100111",
"100001101101100100000101",
"100001101101000000100101",
"100001101100011101000110",
"100001101011111001101000",
"100001101011010110001011",
"100001101010110010101111",
"100001101010001111010100",
"100001101001101011111011",
"100001101001001000100011",
"100001101000100101001100",
"100001101000000001110110",
"100001100111011110100001",
"100001100110111011001101",
"100001100110010111111011",
"100001100101110100101010",
"100001100101010001011001",
"100001100100101110001010",
"100001100100001010111101",
"100001100011100111110000",
"100001100011000100100100",
"100001100010100001011010",
"100001100001111110010001",
"100001100001011011001001",
"100001100000111000000010",
"100001100000010100111100",
"100001011111110001111000",
"100001011111001110110100",
"100001011110101011110010",
"100001011110001000110001",
"100001011101100101110001",
"100001011101000010110010",
"100001011100011111110100",
"100001011011111100110111",
"100001011011011001111100",
"100001011010110111000010",
"100001011010010100001000",
"100001011001110001010000",
"100001011001001110011001",
"100001011000101011100100",
"100001011000001000101111",
"100001010111100101111100",
"100001010111000011001001",
"100001010110100000011000",
"100001010101111101101000",
"100001010101011010111001",
"100001010100111000001011",
"100001010100010101011110",
"100001010011110010110011",
"100001010011010000001000",
"100001010010101101011111",
"100001010010001010110111",
"100001010001101000010000",
"100001010001000101101010",
"100001010000100011000101",
"100001010000000000100001",
"100001001111011101111111",
"100001001110111011011101",
"100001001110011000111101",
"100001001101110110011110",
"100001001101010100000000",
"100001001100110001100011",
"100001001100001111000111",
"100001001011101100101100",
"100001001011001010010010",
"100001001010100111111010",
"100001001010000101100010",
"100001001001100011001100",
"100001001001000000110111",
"100001001000011110100011",
"100001000111111100010000",
"100001000111011001111110",
"100001000110110111101101",
"100001000110010101011110",
"100001000101110011001111",
"100001000101010001000010",
"100001000100101110110101",
"100001000100001100101010",
"100001000011101010100000",
"100001000011001000010111",
"100001000010100110001111",
"100001000010000100001000",
"100001000001100010000011",
"100001000000111111111110",
"100001000000011101111010",
"100000111111111011111000",
"100000111111011001110111",
"100000111110110111110110",
"100000111110010101110111",
"100000111101110011111001",
"100000111101010001111100",
"100000111100110000000001",
"100000111100001110000110",
"100000111011101100001100",
"100000111011001010010100",
"100000111010101000011100",
"100000111010000110100110",
"100000111001100100110000",
"100000111001000010111100",
"100000111000100001001001",
"100000110111111111010111",
"100000110111011101100110",
"100000110110111011110110",
"100000110110011010000111",
"100000110101111000011010",
"100000110101010110101101",
"100000110100110101000001",
"100000110100010011010111",
"100000110011110001101101",
"100000110011010000000101",
"100000110010101110011110",
"100000110010001100111000",
"100000110001101011010011",
"100000110001001001101111",
"100000110000101000001100",
"100000110000000110101010",
"100000101111100101001001",
"100000101111000011101001",
"100000101110100010001011",
"100000101110000000101101",
"100000101101011111010000",
"100000101100111101110101",
"100000101100011100011011",
"100000101011111011000001",
"100000101011011001101001",
"100000101010111000010010",
"100000101010010110111100",
"100000101001110101100111",
"100000101001010100010011",
"100000101000110011000000",
"100000101000010001101110",
"100000100111110000011101",
"100000100111001111001101",
"100000100110101101111111",
"100000100110001100110001",
"100000100101101011100100",
"100000100101001010011001",
"100000100100101001001110",
"100000100100001000000101",
"100000100011100110111101",
"100000100011000101110101",
"100000100010100100101111",
"100000100010000011101010",
"100000100001100010100110",
"100000100001000001100011",
"100000100000100000100001",
"100000011111111111100000",
"100000011111011110100000",
"100000011110111101100001",
"100000011110011100100011",
"100000011101111011100110",
"100000011101011010101010",
"100000011100111001101111",
"100000011100011000110110",
"100000011011110111111101",
"100000011011010111000101",
"100000011010110110001111",
"100000011010010101011001",
"100000011001110100100101",
"100000011001010011110001",
"100000011000110010111111",
"100000011000010010001110",
"100000010111110001011101",
"100000010111010000101110",
"100000010110110000000000",
"100000010110001111010011",
"100000010101101110100110",
"100000010101001101111011",
"100000010100101101010001",
"100000010100001100101000",
"100000010011101100000000",
"100000010011001011011001",
"100000010010101010110011",
"100000010010001010001110",
"100000010001101001101010",
"100000010001001001000111",
"100000010000101000100101",
"100000010000001000000100",
"100000001111100111100100",
"100000001111000111000101",
"100000001110100110100111",
"100000001110000110001011",
"100000001101100101101111",
"100000001101000101010100",
"100000001100100100111010",
"100000001100000100100010",
"100000001011100100001010",
"100000001011000011110011",
"100000001010100011011110",
"100000001010000011001001",
"100000001001100010110101",
"100000001001000010100011",
"100000001000100010010001",
"100000001000000010000001",
"100000000111100001110001",
"100000000111000001100010",
"100000000110100001010101",
"100000000110000001001000",
"100000000101100000111101",
"100000000101000000110010",
"100000000100100000101001",
"100000000100000000100000",
"100000000011100000011001",
"100000000011000000010010",
"100000000010100000001101",
"100000000010000000001000",
"100000000001100000000101",
"100000000001000000000010",
"100000000000100000000001",
"100000000000000000000000"
);

end package fdiv_table;
