library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;


entity PROM is

  port (
    clka  : in  std_logic;
--    wea   : in  std_logic_vector(0 downto 0);
    addra : in  std_logic_vector(6 downto 0);
--    dina  : in  std_logic_vector(31 downto 0);
    douta : out std_logic_vector(31 downto 0));

end PROM;

architecture R_rom of PROM is
--ans(%r1) = 9169
type rom_type is array (0 to 83) of std_logic_vector(31 downto 0);
  constant rom : rom_type:=(
	-- entry:
"11001000000111100000000000000000",	-- 1: 	lli	%sp, 0
"10100100000111110000000000001101",	-- 2: 	addi	%ra, %r0, halt
"11001000000111011100001101010000",	-- 3: 	lli	%hp, 50000
"11001000000000010000000000000011",	-- 4: 	lli	%r1, 3
"11001000000000100000000000000011",	-- 5: 	lli	%r2, 3
"11001000000000110000000000000000",	-- 6: 	lli	%r3, 0
"11001000000001000000000000000000",	-- 7: 	lli	%r4, 0
"00111111111111100000000000000000",	-- 8: 	sw	%ra, [%sp + 0]
"10100111110111100000000000000001",	-- 9: 	addi	%sp, %sp, 1
"01011000000000000000000000001110",	-- 10: 	jal	f.46
"10101011110111100000000000000001",	-- 11: 	subi	%sp, %sp, 1
"00111011110111110000000000000000",	-- 12: 	lw	%ra, [%sp + 0]
"01010100000000000000000001010100",	-- 13: 	j	yj_print_int
	-- halt:
"11000000000000000000000000000000",	-- 14: 	halt
	-- f.46:
"11001000000001010000000001100100",	-- 15: 	lli	%r5, 100
"00110000011001010000000000100111",	-- 16: 	bgt	%r3, %r5, bgt_else.97
"11001000000001010010011100010000",	-- 17: 	lli	%r5, 10000
"00110000010001010000000000011110",	-- 18: 	bgt	%r2, %r5, bgt_else.98
"11001000000001010010011100010000",	-- 19: 	lli	%r5, 10000
"00110000001001010000000000010010",	-- 20: 	bgt	%r1, %r5, bgt_else.99
"00110000010000010000000000001001",	-- 21: 	bgt	%r2, %r1, bgt_else.100
"10001100001000100010100000000000",	-- 22: 	mul	%r5, %r1, %r2
"10000100010000010001000000000000",	-- 23: 	add	%r2, %r2, %r1
"11001000000000010000000000000001",	-- 24: 	lli	%r1, 1
"10000100011000010001100000000000",	-- 25: 	add	%r3, %r3, %r1
"11001000000000010000000000000001",	-- 26: 	lli	%r1, 1
"10001000100000010010000000000000",	-- 27: 	sub	%r4, %r4, %r1
"10000100000001010000100000000000",	-- 28: 	add	%r1, %r0, %r5
"01010100000000000000000000001110",	-- 29: 	j	f.46
	-- bgt_else.100:
"10001100001000100010100000000000",	-- 30: 	mul	%r5, %r1, %r2
"10001000010000010001000000000000",	-- 31: 	sub	%r2, %r2, %r1
"11001000000000010000000000000001",	-- 32: 	lli	%r1, 1
"10000100011000010001100000000000",	-- 33: 	add	%r3, %r3, %r1
"11001000000000010000000000000001",	-- 34: 	lli	%r1, 1
"10001000100000010010000000000000",	-- 35: 	sub	%r4, %r4, %r1
"10000100000001010000100000000000",	-- 36: 	add	%r1, %r0, %r5
"01010100000000000000000000001110",	-- 37: 	j	f.46
	-- bgt_else.99:
"10001100001000100001000000000000",	-- 38: 	mul	%r2, %r1, %r2
"01000000001000010000000000000001",	-- 39: 	sra	%r1, %r1, 1
"11001000000001010000000000000001",	-- 40: 	lli	%r5, 1
"10000100011001010001100000000000",	-- 41: 	add	%r3, %r3, %r5
"11001000000001010000000000000001",	-- 42: 	lli	%r5, 1
"10001000100001010010000000000000",	-- 43: 	sub	%r4, %r4, %r5
"10000100000000101101000000000000",	-- 44: 	add	%r26, %r0, %r2
"10000100000000010001000000000000",	-- 45: 	add	%r2, %r0, %r1
"10000100000110100000100000000000",	-- 46: 	add	%r1, %r0, %r26
"01010100000000000000000000001110",	-- 47: 	j	f.46
	-- bgt_else.98:
"10001100001000100000100000000000",	-- 48: 	mul	%r1, %r1, %r2
"01000000010000100000000000000001",	-- 49: 	sra	%r2, %r2, 1
"11001000000001010000000000000001",	-- 50: 	lli	%r5, 1
"10000100011001010001100000000000",	-- 51: 	add	%r3, %r3, %r5
"11001000000001010000000000000001",	-- 52: 	lli	%r5, 1
"10001000100001010010000000000000",	-- 53: 	sub	%r4, %r4, %r5
"01010100000000000000000000001110",	-- 54: 	j	f.46
	-- bgt_else.97:
"11001000000001010000000001100101",	-- 55: 	lli	%r5, 101
"00110000011001010000000000011010",	-- 56: 	bgt	%r3, %r5, bgt_else.101
"11001000000001011111111110011100",	-- 57: 	lli	%r5, -100
"11001100000001011111111111111111",	-- 58: 	lhi	%r5, -100
"00110000101001000000000000000100",	-- 59: 	bgt	%r5, %r4, bgt_else.102
"11001000000000011111111111111100",	-- 60: 	lli	%r1, -4
"11001100000000011111111111111111",	-- 61: 	lhi	%r1, -4
"01001111111000000000000000000000",	-- 62: 	jr	%ra
	-- bgt_else.102:
"11001000000001011111111110011011",	-- 63: 	lli	%r5, -101
"11001100000001011111111111111111",	-- 64: 	lhi	%r5, -101
"00110000101001000000000000001110",	-- 65: 	bgt	%r5, %r4, bgt_else.103
"11001000000001010000000001100101",	-- 66: 	lli	%r5, 101
"00101000011001010000000000001001",	-- 67: 	bneq	%r3, %r5, bneq_else.104
"11001000000000111111111110011011",	-- 68: 	lli	%r3, -101
"11001100000000111111111111111111",	-- 69: 	lhi	%r3, -101
"00101000100000110000000000000011",	-- 70: 	bneq	%r4, %r3, bneq_else.105
"10000100001000100000100000000000",	-- 71: 	add	%r1, %r1, %r2
"01001111111000000000000000000000",	-- 72: 	jr	%ra
	-- bneq_else.105:
"11001000000000011111111111111111",	-- 73: 	lli	%r1, -1
"11001100000000011111111111111111",	-- 74: 	lhi	%r1, -1
"01001111111000000000000000000000",	-- 75: 	jr	%ra
	-- bneq_else.104:
"11001000000000011111111111111110",	-- 76: 	lli	%r1, -2
"11001100000000011111111111111111",	-- 77: 	lhi	%r1, -2
"01001111111000000000000000000000",	-- 78: 	jr	%ra
	-- bgt_else.103:
"11001000000000011111111111111101",	-- 79: 	lli	%r1, -3
"11001100000000011111111111111111",	-- 80: 	lhi	%r1, -3
"01001111111000000000000000000000",	-- 81: 	jr	%ra
	-- bgt_else.101:
"11001000000000011111111111111011",	-- 82: 	lli	%r1, -5
"11001100000000011111111111111111",	-- 83: 	lhi	%r1, -5
"01001111111000000000000000000000"	-- 84: 	jr	%ra
);

signal shortened : std_logic_vector(6 downto 0):=(others=>'0');
begin  -- R_rom
  shortened<=addra(6 downto 0);
    douta<=rom(conv_integer(shortened));
end R_rom;
